VERSION 5.8 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

PROPERTYDEFINITIONS
  MACRO expanded_util REAL ;
  MACRO previous_effective_target_usage REAL ;
END PROPERTYDEFINITIONS

LAYER NWELL
  TYPE MASTERSLICE ;
END NWELL

LAYER LVTIMP
  TYPE IMPLANT ;
END LVTIMP

LAYER PO
  TYPE MASTERSLICE ;
END PO

LAYER M1
  TYPE ROUTING ;
  MASK 2 ;
  DIRECTION VERTICAL ;
  PITCH 0.074 ;
  WIDTH 0.034 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.034 WRONGDIRECTION ;" ;
END M1

LAYER VIA1
  TYPE CUT ;
END VIA1

LAYER M2
  TYPE ROUTING ;
  MASK 2 ;
  DIRECTION HORIZONTAL ;
  PITCH 0.06 ;
  WIDTH 0.034 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.034 WRONGDIRECTION ;" ;
END M2

LAYER VIA2
  TYPE CUT ;
END VIA2

LAYER M3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.074 ;
  WIDTH 0.034 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.034 WRONGDIRECTION ;" ;
END M3

LAYER VIA3
  TYPE CUT ;
END VIA3

LAYER M4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.074 ;
  WIDTH 0.06 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.06 WRONGDIRECTION ;" ;
END M4

LAYER VIA4
  TYPE CUT ;
END VIA4

LAYER M5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.12 ;
  WIDTH 0.06 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.06 WRONGDIRECTION ;" ;
END M5

LAYER VIA5
  TYPE CUT ;
END VIA5

LAYER M6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.12 ;
  WIDTH 0.06 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.06 WRONGDIRECTION ;" ;
END M6

LAYER VIA6
  TYPE CUT ;
END VIA6

LAYER M7
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.12 ;
  WIDTH 0.06 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.06 WRONGDIRECTION ;" ;
END M7

LAYER VIA7
  TYPE CUT ;
END VIA7

LAYER M8
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.12 ;
  WIDTH 0.06 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.06 WRONGDIRECTION ;" ;
END M8

LAYER VIA8
  TYPE CUT ;
END VIA8

LAYER M9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.12 ;
  WIDTH 0.06 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.06 WRONGDIRECTION ;" ;
END M9

LAYER VIARDL
  TYPE CUT ;
END VIARDL

LAYER MRDL
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.6 ;
  WIDTH 2 ;
  PROPERTY LEF58_WIDTH "WIDTH 2 WRONGDIRECTION ;" ;
END MRDL

LAYER DIFF
  TYPE MASTERSLICE ;
END DIFF

LAYER FIN
  TYPE MASTERSLICE ;
END FIN

LAYER DNW
  TYPE MASTERSLICE ;
END DNW

LAYER PIMP
  TYPE MASTERSLICE ;
END PIMP

LAYER NIMP
  TYPE MASTERSLICE ;
END NIMP

LAYER DIFF_15
  TYPE MASTERSLICE ;
END DIFF_15

LAYER PAD
  TYPE MASTERSLICE ;
END PAD

LAYER ESD
  TYPE MASTERSLICE ;
END ESD

LAYER SBLK
  TYPE MASTERSLICE ;
END SBLK

LAYER CPO
  TYPE MASTERSLICE ;
END CPO

LAYER CTM1
  TYPE MASTERSLICE ;
END CTM1

LAYER VIA0
  TYPE MASTERSLICE ;
END VIA0

LAYER HVTIMP
  TYPE IMPLANT ;
END HVTIMP

LAYER M1PIN
  TYPE MASTERSLICE ;
END M1PIN

LAYER M2PIN
  TYPE MASTERSLICE ;
END M2PIN

LAYER M3PIN
  TYPE MASTERSLICE ;
END M3PIN

LAYER M4PIN
  TYPE MASTERSLICE ;
END M4PIN

LAYER M5PIN
  TYPE MASTERSLICE ;
END M5PIN

LAYER M6PIN
  TYPE MASTERSLICE ;
END M6PIN

LAYER M7PIN
  TYPE MASTERSLICE ;
END M7PIN

LAYER M8PIN
  TYPE MASTERSLICE ;
END M8PIN

LAYER M9PIN
  TYPE MASTERSLICE ;
END M9PIN

LAYER MRPIN
  TYPE MASTERSLICE ;
END MRPIN

LAYER HOTNWL
  TYPE MASTERSLICE ;
END HOTNWL

LAYER DIOD
  TYPE MASTERSLICE ;
END DIOD

LAYER BJTDMY
  TYPE MASTERSLICE ;
END BJTDMY

LAYER RNW
  TYPE MASTERSLICE ;
END RNW

LAYER RMARK
  TYPE MASTERSLICE ;
END RMARK

LAYER prBoundary
  TYPE MASTERSLICE ;
END prBoundary

LAYER LOGO
  TYPE MASTERSLICE ;
END LOGO

LAYER IP
  TYPE MASTERSLICE ;
END IP

LAYER RM1
  TYPE MASTERSLICE ;
END RM1

LAYER RM2
  TYPE MASTERSLICE ;
END RM2

LAYER RM3
  TYPE MASTERSLICE ;
END RM3

LAYER RM4
  TYPE MASTERSLICE ;
END RM4

LAYER RM5
  TYPE MASTERSLICE ;
END RM5

LAYER RM6
  TYPE MASTERSLICE ;
END RM6

LAYER RM7
  TYPE MASTERSLICE ;
END RM7

LAYER RM8
  TYPE MASTERSLICE ;
END RM8

LAYER RM9
  TYPE MASTERSLICE ;
END RM9

LAYER DIFF_25
  TYPE MASTERSLICE ;
END DIFF_25

VIA VIA12SQ_C
  LAYER M1 ;
    RECT -0.055 -0.017 0.055 0.017 ;
  LAYER VIA1 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M2 ;
    RECT -0.017 -0.055 0.017 0.055 ;
END VIA12SQ_C

VIA VIA12BAR1_C
  LAYER M1 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA1 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER M2 ;
    RECT -0.017 -0.075 0.017 0.075 ;
END VIA12BAR1_C

VIA VIA12BAR2_C
  LAYER M1 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA1 ;
    RECT -0.03 -0.015 0.03 0.015 ;
  LAYER M2 ;
    RECT -0.032 -0.04 0.032 0.04 ;
END VIA12BAR2_C

VIA VIA12LG_C
  LAYER M1 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA1 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA12LG_C

VIA VIA12SQ
  LAYER M1 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA1 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
END VIA12SQ

VIA VIA12BAR1
  LAYER M1 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA1 ;
    RECT -0.03 -0.015 0.03 0.015 ;
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
END VIA12BAR1

VIA VIA12BAR2
  LAYER M1 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA1 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA12BAR2

VIA VIA12LG
  LAYER M1 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA1 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA12LG

VIA VIA1_32SQ_C
  LAYER M1 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA1 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M2 ;
    RECT -0.017 -0.075 0.017 0.075 ;
END VIA1_32SQ_C

VIA VIA1_32BAR1_C
  LAYER M1 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA1 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER M2 ;
    RECT -0.017 -0.075 0.017 0.075 ;
END VIA1_32BAR1_C

VIA VIA1_32BAR2_C
  LAYER M1 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA1 ;
    RECT -0.03 -0.015 0.03 0.015 ;
  LAYER M2 ;
    RECT -0.032 -0.04 0.032 0.04 ;
END VIA1_32BAR2_C

VIA VIA1_32LG_C
  LAYER M1 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA1 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA1_32LG_C

VIA VIA1_32SQ
  LAYER M1 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA1 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
END VIA1_32SQ

VIA VIA1_32BAR1
  LAYER M1 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA1 ;
    RECT -0.03 -0.015 0.03 0.015 ;
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
END VIA1_32BAR1

VIA VIA1_32BAR2
  LAYER M1 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA1 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA1_32BAR2

VIA VIA1_32LG
  LAYER M1 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA1 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA1_32LG

VIA VIA12_3SQ_C
  LAYER M1 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA1 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M2 ;
    RECT -0.017 -0.075 0.017 0.075 ;
END VIA12_3SQ_C

VIA VIA12_3BAR1_C
  LAYER M1 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA1 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER M2 ;
    RECT -0.017 -0.075 0.017 0.075 ;
END VIA12_3BAR1_C

VIA VIA12_3BAR2_C
  LAYER M1 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA1 ;
    RECT -0.03 -0.015 0.03 0.015 ;
  LAYER M2 ;
    RECT -0.032 -0.04 0.032 0.04 ;
END VIA12_3BAR2_C

VIA VIA12_3LG_C
  LAYER M1 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA1 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA12_3LG_C

VIA VIA12_3SQ
  LAYER M1 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA1 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
END VIA12_3SQ

VIA VIA12_3BAR1
  LAYER M1 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA1 ;
    RECT -0.03 -0.015 0.03 0.015 ;
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
END VIA12_3BAR1

VIA VIA12_3BAR2
  LAYER M1 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA1 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA12_3BAR2

VIA VIA12_3LG
  LAYER M1 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA1 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA12_3LG

VIA VIA1_32_3SQ_C
  LAYER M1 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA1 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M2 ;
    RECT -0.017 -0.075 0.017 0.075 ;
END VIA1_32_3SQ_C

VIA VIA1_32_3BAR1_C
  LAYER M1 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA1 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER M2 ;
    RECT -0.017 -0.075 0.017 0.075 ;
END VIA1_32_3BAR1_C

VIA VIA1_32_3BAR2_C
  LAYER M1 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA1 ;
    RECT -0.03 -0.015 0.03 0.015 ;
  LAYER M2 ;
    RECT -0.032 -0.04 0.032 0.04 ;
END VIA1_32_3BAR2_C

VIA VIA1_32_3LG_C
  LAYER M1 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA1 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA1_32_3LG_C

VIA VIA1_32_3SQ
  LAYER M1 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA1 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
END VIA1_32_3SQ

VIA VIA1_32_3BAR1
  LAYER M1 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA1 ;
    RECT -0.03 -0.015 0.03 0.015 ;
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
END VIA1_32_3BAR1

VIA VIA1_32_3BAR2
  LAYER M1 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA1 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA1_32_3BAR2

VIA VIA1_32_3LG
  LAYER M1 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA1 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA1_32_3LG

VIA VIA23SQ_C
  LAYER M2 ;
    RECT -0.055 -0.017 0.055 0.017 ;
  LAYER VIA2 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M3 ;
    RECT -0.017 -0.055 0.017 0.055 ;
END VIA23SQ_C

VIA VIA23BAR1_C
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA2 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER M3 ;
    RECT -0.017 -0.075 0.017 0.075 ;
END VIA23BAR1_C

VIA VIA23BAR2_C
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA2 ;
    RECT -0.03 -0.015 0.03 0.015 ;
  LAYER M3 ;
    RECT -0.032 -0.04 0.032 0.04 ;
END VIA23BAR2_C

VIA VIA23LG_C
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA2 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M3 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA23LG_C

VIA VIA23SQ
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA2 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M3 ;
    RECT -0.075 -0.017 0.075 0.017 ;
END VIA23SQ

VIA VIA23BAR1
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA2 ;
    RECT -0.03 -0.015 0.03 0.015 ;
  LAYER M3 ;
    RECT -0.075 -0.017 0.075 0.017 ;
END VIA23BAR1

VIA VIA23BAR2
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA2 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER M3 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA23BAR2

VIA VIA23LG
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA2 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M3 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA23LG

VIA VIA2_33SQ_C
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA2 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M3 ;
    RECT -0.017 -0.075 0.017 0.075 ;
END VIA2_33SQ_C

VIA VIA2_33BAR1_C
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA2 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER M3 ;
    RECT -0.017 -0.075 0.017 0.075 ;
END VIA2_33BAR1_C

VIA VIA2_33BAR2_C
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA2 ;
    RECT -0.03 -0.015 0.03 0.015 ;
  LAYER M3 ;
    RECT -0.032 -0.04 0.032 0.04 ;
END VIA2_33BAR2_C

VIA VIA2_33LG_C
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA2 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M3 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA2_33LG_C

VIA VIA2_33SQ
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA2 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M3 ;
    RECT -0.075 -0.017 0.075 0.017 ;
END VIA2_33SQ

VIA VIA2_33BAR1
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA2 ;
    RECT -0.03 -0.015 0.03 0.015 ;
  LAYER M3 ;
    RECT -0.075 -0.017 0.075 0.017 ;
END VIA2_33BAR1

VIA VIA2_33BAR2
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA2 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER M3 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA2_33BAR2

VIA VIA2_33LG
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA2 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M3 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA2_33LG

VIA VIA23_3SQ_C
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA2 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M3 ;
    RECT -0.017 -0.075 0.017 0.075 ;
END VIA23_3SQ_C

VIA VIA23_3BAR1_C
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA2 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER M3 ;
    RECT -0.017 -0.075 0.017 0.075 ;
END VIA23_3BAR1_C

VIA VIA23_3BAR2_C
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA2 ;
    RECT -0.03 -0.015 0.03 0.015 ;
  LAYER M3 ;
    RECT -0.032 -0.04 0.032 0.04 ;
END VIA23_3BAR2_C

VIA VIA23_3LG_C
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA2 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M3 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA23_3LG_C

VIA VIA23_3SQ
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA2 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M3 ;
    RECT -0.075 -0.017 0.075 0.017 ;
END VIA23_3SQ

VIA VIA23_3BAR1
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA2 ;
    RECT -0.03 -0.015 0.03 0.015 ;
  LAYER M3 ;
    RECT -0.075 -0.017 0.075 0.017 ;
END VIA23_3BAR1

VIA VIA23_3BAR2
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA2 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER M3 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA23_3BAR2

VIA VIA23_3LG
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA2 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M3 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA23_3LG

VIA VIA2_33_3SQ_C
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA2 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M3 ;
    RECT -0.017 -0.075 0.017 0.075 ;
END VIA2_33_3SQ_C

VIA VIA2_33_3BAR1_C
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA2 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER M3 ;
    RECT -0.017 -0.075 0.017 0.075 ;
END VIA2_33_3BAR1_C

VIA VIA2_33_3BAR2_C
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA2 ;
    RECT -0.03 -0.015 0.03 0.015 ;
  LAYER M3 ;
    RECT -0.032 -0.04 0.032 0.04 ;
END VIA2_33_3BAR2_C

VIA VIA2_33_3LG_C
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA2 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M3 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA2_33_3LG_C

VIA VIA2_33_3SQ
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA2 ;
    RECT -0.015 -0.015 0.015 0.015 ;
  LAYER M3 ;
    RECT -0.075 -0.017 0.075 0.017 ;
END VIA2_33_3SQ

VIA VIA2_33_3BAR1
  LAYER M2 ;
    RECT -0.075 -0.017 0.075 0.017 ;
  LAYER VIA2 ;
    RECT -0.03 -0.015 0.03 0.015 ;
  LAYER M3 ;
    RECT -0.075 -0.017 0.075 0.017 ;
END VIA2_33_3BAR1

VIA VIA2_33_3BAR2
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA2 ;
    RECT -0.015 -0.03 0.015 0.03 ;
  LAYER M3 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA2_33_3BAR2

VIA VIA2_33_3LG
  LAYER M2 ;
    RECT -0.04 -0.032 0.04 0.032 ;
  LAYER VIA2 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M3 ;
    RECT -0.04 -0.032 0.04 0.032 ;
END VIA2_33_3LG

VIA VIA34SQ_C
  LAYER M3 ;
    RECT -0.037 -0.035 0.037 0.035 ;
  LAYER VIA3 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M4 ;
    RECT -0.035 -0.037 0.035 0.037 ;
END VIA34SQ_C

VIA VIA34BAR1_C
  LAYER M3 ;
    RECT -0.065 -0.035 0.065 0.035 ;
  LAYER VIA3 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER M4 ;
    RECT -0.065 -0.035 0.065 0.035 ;
END VIA34BAR1_C

VIA VIA34BAR2_C
  LAYER M3 ;
    RECT -0.035 -0.065 0.035 0.065 ;
  LAYER VIA3 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER M4 ;
    RECT -0.035 -0.065 0.035 0.065 ;
END VIA34BAR2_C

VIA VIA34LG_C
  LAYER M3 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER VIA3 ;
    RECT -0.06 -0.06 0.06 0.06 ;
  LAYER M4 ;
    RECT -0.065 -0.065 0.065 0.065 ;
END VIA34LG_C

VIA VIA34SQ
  LAYER M3 ;
    RECT -0.037 -0.035 0.037 0.035 ;
  LAYER VIA3 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M4 ;
    RECT -0.037 -0.035 0.037 0.035 ;
END VIA34SQ

VIA VIA34BAR1
  LAYER M3 ;
    RECT -0.065 -0.035 0.065 0.035 ;
  LAYER VIA3 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER M4 ;
    RECT -0.065 -0.035 0.065 0.035 ;
END VIA34BAR1

VIA VIA34BAR2
  LAYER M3 ;
    RECT -0.035 -0.065 0.035 0.065 ;
  LAYER VIA3 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER M4 ;
    RECT -0.035 -0.065 0.035 0.065 ;
END VIA34BAR2

VIA VIA34LG
  LAYER M3 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER VIA3 ;
    RECT -0.06 -0.06 0.06 0.06 ;
  LAYER M4 ;
    RECT -0.065 -0.065 0.065 0.065 ;
END VIA34LG

VIA VIA3_34SQ_C
  LAYER M3 ;
    RECT -0.037 -0.035 0.037 0.035 ;
  LAYER VIA3 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M4 ;
    RECT -0.035 -0.037 0.035 0.037 ;
END VIA3_34SQ_C

VIA VIA3_34BAR1_C
  LAYER M3 ;
    RECT -0.065 -0.035 0.065 0.035 ;
  LAYER VIA3 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER M4 ;
    RECT -0.065 -0.035 0.065 0.035 ;
END VIA3_34BAR1_C

VIA VIA3_34BAR2_C
  LAYER M3 ;
    RECT -0.035 -0.065 0.035 0.065 ;
  LAYER VIA3 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER M4 ;
    RECT -0.035 -0.065 0.035 0.065 ;
END VIA3_34BAR2_C

VIA VIA3_34LG_C
  LAYER M3 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER VIA3 ;
    RECT -0.06 -0.06 0.06 0.06 ;
  LAYER M4 ;
    RECT -0.065 -0.065 0.065 0.065 ;
END VIA3_34LG_C

VIA VIA3_34SQ
  LAYER M3 ;
    RECT -0.037 -0.035 0.037 0.035 ;
  LAYER VIA3 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M4 ;
    RECT -0.037 -0.035 0.037 0.035 ;
END VIA3_34SQ

VIA VIA3_34BAR1
  LAYER M3 ;
    RECT -0.065 -0.035 0.065 0.035 ;
  LAYER VIA3 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER M4 ;
    RECT -0.065 -0.035 0.065 0.035 ;
END VIA3_34BAR1

VIA VIA3_34BAR2
  LAYER M3 ;
    RECT -0.035 -0.065 0.035 0.065 ;
  LAYER VIA3 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER M4 ;
    RECT -0.035 -0.065 0.035 0.065 ;
END VIA3_34BAR2

VIA VIA3_4LG
  LAYER M3 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER VIA3 ;
    RECT -0.06 -0.06 0.06 0.06 ;
  LAYER M4 ;
    RECT -0.065 -0.065 0.065 0.065 ;
END VIA3_4LG

VIA VIA45BAR1_C
  LAYER M4 ;
    RECT -0.065 -0.035 0.065 0.035 ;
  LAYER VIA4 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER M5 ;
    RECT -0.065 -0.035 0.065 0.035 ;
END VIA45BAR1_C

VIA VIA45BAR2_C
  LAYER M4 ;
    RECT -0.035 -0.065 0.035 0.065 ;
  LAYER VIA4 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER M5 ;
    RECT -0.035 -0.065 0.035 0.065 ;
END VIA45BAR2_C

VIA VIA45LG_C
  LAYER M4 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER VIA4 ;
    RECT -0.06 -0.06 0.06 0.06 ;
  LAYER M5 ;
    RECT -0.065 -0.065 0.065 0.065 ;
END VIA45LG_C

VIA VIA45SQ
  LAYER M4 ;
    RECT -0.037 -0.035 0.037 0.035 ;
  LAYER VIA4 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M5 ;
    RECT -0.037 -0.035 0.037 0.035 ;
END VIA45SQ

VIA VIA45BAR1
  LAYER M4 ;
    RECT -0.065 -0.035 0.065 0.035 ;
  LAYER VIA4 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER M5 ;
    RECT -0.065 -0.035 0.065 0.035 ;
END VIA45BAR1

VIA VIA45BAR2
  LAYER M4 ;
    RECT -0.035 -0.065 0.035 0.065 ;
  LAYER VIA4 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER M5 ;
    RECT -0.035 -0.065 0.035 0.065 ;
END VIA45BAR2

VIA VIA45LG
  LAYER M4 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER VIA4 ;
    RECT -0.06 -0.06 0.06 0.06 ;
  LAYER M5 ;
    RECT -0.065 -0.065 0.065 0.065 ;
END VIA45LG

VIA VIA56SQ_C
  LAYER M5 ;
    RECT -0.037 -0.035 0.037 0.035 ;
  LAYER VIA5 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M6 ;
    RECT -0.035 -0.037 0.035 0.037 ;
END VIA56SQ_C

VIA VIA56BAR1_C
  LAYER M5 ;
    RECT -0.065 -0.035 0.065 0.035 ;
  LAYER VIA5 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER M6 ;
    RECT -0.065 -0.035 0.065 0.035 ;
END VIA56BAR1_C

VIA VIA56BAR2_C
  LAYER M5 ;
    RECT -0.035 -0.065 0.035 0.065 ;
  LAYER VIA5 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER M6 ;
    RECT -0.035 -0.065 0.035 0.065 ;
END VIA56BAR2_C

VIA VIA56LG_C
  LAYER M5 ;
    RECT -0.035 -0.065 0.035 0.065 ;
  LAYER VIA5 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER M6 ;
    RECT -0.035 -0.065 0.035 0.065 ;
END VIA56LG_C

VIA VIA56SQ
  LAYER M5 ;
    RECT -0.035 -0.035 0.035 0.035 ;
  LAYER VIA5 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M6 ;
    RECT -0.035 -0.035 0.035 0.035 ;
END VIA56SQ

VIA VIA56BAR1
  LAYER M5 ;
    RECT -0.065 -0.035 0.065 0.035 ;
  LAYER VIA5 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER M6 ;
    RECT -0.065 -0.035 0.065 0.035 ;
END VIA56BAR1

VIA VIA56BAR2
  LAYER M5 ;
    RECT -0.035 -0.065 0.035 0.065 ;
  LAYER VIA5 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER M6 ;
    RECT -0.035 -0.065 0.035 0.065 ;
END VIA56BAR2

VIA VIA56LG
  LAYER M5 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER VIA5 ;
    RECT -0.06 -0.06 0.06 0.06 ;
  LAYER M6 ;
    RECT -0.065 -0.065 0.065 0.065 ;
END VIA56LG

VIA VIA67SQ_C
  LAYER M6 ;
    RECT -0.037 -0.035 0.037 0.035 ;
  LAYER VIA6 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M7 ;
    RECT -0.035 -0.037 0.035 0.037 ;
END VIA67SQ_C

VIA VIA67BAR1_C
  LAYER M6 ;
    RECT -0.065 -0.035 0.065 0.035 ;
  LAYER VIA6 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER M7 ;
    RECT -0.065 -0.035 0.065 0.035 ;
END VIA67BAR1_C

VIA VIA67SQ
  LAYER M6 ;
    RECT -0.037 -0.035 0.037 0.035 ;
  LAYER VIA6 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M7 ;
    RECT -0.037 -0.035 0.037 0.035 ;
END VIA67SQ

VIA VIA67BAR1
  LAYER M6 ;
    RECT -0.065 -0.035 0.065 0.035 ;
  LAYER VIA6 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER M7 ;
    RECT -0.065 -0.035 0.065 0.035 ;
END VIA67BAR1

VIA VIA67BAR2
  LAYER M6 ;
    RECT -0.035 -0.065 0.035 0.065 ;
  LAYER VIA6 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER M7 ;
    RECT -0.035 -0.065 0.035 0.065 ;
END VIA67BAR2

VIA VIA67LG
  LAYER M6 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER VIA6 ;
    RECT -0.06 -0.06 0.06 0.06 ;
  LAYER M7 ;
    RECT -0.065 -0.065 0.065 0.065 ;
END VIA67LG

VIA VIA78SQ_C
  LAYER M7 ;
    RECT -0.037 -0.035 0.037 0.035 ;
  LAYER VIA7 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M8 ;
    RECT -0.035 -0.037 0.035 0.037 ;
END VIA78SQ_C

VIA VIA78BAR1_C
  LAYER M7 ;
    RECT -0.065 -0.035 0.065 0.035 ;
  LAYER VIA7 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER M8 ;
    RECT -0.065 -0.035 0.065 0.035 ;
END VIA78BAR1_C

VIA VIA78BAR2_C
  LAYER M7 ;
    RECT -0.037 -0.067 0.037 0.067 ;
  LAYER VIA7 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER M8 ;
    RECT -0.037 -0.067 0.037 0.067 ;
END VIA78BAR2_C

VIA VIA78LG_C
  LAYER M7 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER VIA7 ;
    RECT -0.06 -0.06 0.06 0.06 ;
  LAYER M8 ;
    RECT -0.065 -0.065 0.065 0.065 ;
END VIA78LG_C

VIA VIA78SQ
  LAYER M7 ;
    RECT -0.037 -0.035 0.037 0.035 ;
  LAYER VIA7 ;
    RECT -0.03 -0.03 0.03 0.03 ;
  LAYER M8 ;
    RECT -0.037 -0.035 0.037 0.035 ;
END VIA78SQ

VIA VIA78BAR1
  LAYER M7 ;
    RECT -0.065 -0.035 0.065 0.035 ;
  LAYER VIA7 ;
    RECT -0.06 -0.03 0.06 0.03 ;
  LAYER M8 ;
    RECT -0.065 -0.035 0.065 0.035 ;
END VIA78BAR1

VIA VIA78BAR2
  LAYER M7 ;
    RECT -0.035 -0.065 0.035 0.065 ;
  LAYER VIA7 ;
    RECT -0.03 -0.06 0.03 0.06 ;
  LAYER M8 ;
    RECT -0.035 -0.065 0.035 0.065 ;
END VIA78BAR2

VIA VIA78LG
  LAYER M7 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER VIA7 ;
    RECT -0.06 -0.06 0.06 0.06 ;
  LAYER M8 ;
    RECT -0.065 -0.065 0.065 0.065 ;
END VIA78LG

VIA VIA89_C
  LAYER M8 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER VIA8 ;
    RECT -0.06 -0.06 0.06 0.06 ;
  LAYER M9 ;
    RECT -0.065 -0.065 0.065 0.065 ;
END VIA89_C

VIA VIA89
  LAYER M8 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER VIA8 ;
    RECT -0.06 -0.06 0.06 0.06 ;
  LAYER M9 ;
    RECT -0.065 -0.065 0.065 0.065 ;
END VIA89

VIA VIA9RDL
  LAYER M9 ;
    RECT -1.5 -1.5 1.5 1.5 ;
  LAYER VIARDL ;
    RECT -1 -1 1 1 ;
  LAYER MRDL ;
    RECT -1.5 -1.5 1.5 1.5 ;
END VIA9RDL

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.074 BY 0.6 ;
END unit

MACRO SAEDRVT14_FSDPSYNSBQ_V2LP_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.22 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.17 0.225 0.2 0.255 ;
      LAYER M2 ;
        RECT 0.146 0.223 0.382 0.257 ;
        RECT MASK 1 0.146 0.223 0.382 0.257 ;
    END
  END SD
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 0.176 0.424 0.418 ;
        RECT MASK 1 0.39 0.176 0.424 0.418 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.76 0.263 0.794 0.458 ;
        RECT MASK 1 0.76 0.263 0.794 0.458 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.686 0.224 0.72 0.488 ;
        RECT MASK 1 0.686 0.224 0.72 0.488 ;
    END
  END SE
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.946 0.285 1.976 0.315 ;
      LAYER M2 ;
        RECT 1.861 0.283 2.098 0.317 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 2.092 0.088 2.126 0.488 ;
        RECT 2.092 0.088 2.126 0.488 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 2.262 0.647 ;
        RECT MASK 1 -0.042 0.553 2.262 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 2.262 0.047 ;
        RECT MASK 1 -0.042 -0.047 2.262 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 1.87 0.464 2.022 0.498 ;
      RECT MASK 1 1.87 0.136 1.904 0.464 ;
      RECT MASK 1 1.87 0.102 2 0.136 ;
      RECT MASK 1 0.316 0.464 0.534 0.498 ;
      RECT MASK 1 0.316 0.136 0.35 0.464 ;
      RECT MASK 1 0.222 0.102 0.464 0.136 ;
      RECT MASK 1 0.094 0.464 0.276 0.498 ;
      RECT MASK 1 0.094 0.088 0.128 0.464 ;
      RECT MASK 1 0.242 0.224 0.276 0.464 ;
      RECT MASK 1 1.485 0.462 1.682 0.496 ;
      RECT MASK 1 1.648 0.136 1.682 0.462 ;
      RECT MASK 1 1.426 0.102 1.682 0.136 ;
      RECT MASK 1 1.209 0.462 1.391 0.496 ;
      RECT MASK 1 1.209 0.136 1.243 0.462 ;
      RECT MASK 1 1.209 0.102 1.386 0.136 ;
      RECT MASK 1 1.13 0.395 1.164 0.488 ;
      RECT MASK 1 1.056 0.361 1.164 0.395 ;
      RECT MASK 1 1.056 0.088 1.09 0.361 ;
      RECT MASK 1 0.834 0.088 0.868 0.488 ;
      RECT MASK 1 0.612 0.395 0.646 0.488 ;
      RECT MASK 1 0.538 0.361 0.646 0.395 ;
      RECT MASK 1 0.538 0.088 0.572 0.361 ;
      RECT MASK 1 1.796 0.118 1.83 0.458 ;
      RECT MASK 1 1.722 0.118 1.756 0.458 ;
      RECT MASK 1 0.982 0.224 1.016 0.458 ;
      RECT MASK 1 1.426 0.199 1.46 0.43 ;
      RECT MASK 1 2.018 0.163 2.052 0.418 ;
      RECT MASK 1 1.288 0.263 1.334 0.418 ;
      RECT MASK 1 0.908 0.088 0.942 0.418 ;
      RECT MASK 1 1.944 0.259 1.978 0.413 ;
      RECT MASK 1 1.574 0.199 1.608 0.377 ;
      RECT MASK 1 1.5 0.199 1.534 0.377 ;
      RECT MASK 1 0.464 0.176 0.498 0.37 ;
      RECT MASK 1 0.168 0.171 0.202 0.365 ;
      RECT MASK 1 1.13 0.158 1.164 0.313 ;
      RECT MASK 1 0.612 0.118 0.646 0.313 ;
    LAYER M2 ;
      RECT MASK 1 0.938 0.343 1.942 0.377 ;
      RECT MASK 1 1.08 0.223 1.835 0.257 ;
      RECT MASK 1 0.46 0.223 0.924 0.257 ;
      RECT MASK 1 0.477 0.103 0.966 0.137 ;
    LAYER VIA1 ;
      RECT 1.872 0.345 1.902 0.375 ;
      RECT 1.428 0.345 1.458 0.375 ;
      RECT 0.984 0.345 1.014 0.375 ;
      RECT 1.724 0.285 1.754 0.315 ;
      RECT 1.576 0.285 1.606 0.315 ;
      RECT 1.295 0.285 1.325 0.315 ;
      RECT 1.058 0.285 1.088 0.315 ;
      RECT 1.798 0.225 1.828 0.255 ;
      RECT 1.502 0.225 1.532 0.255 ;
      RECT 1.132 0.225 1.162 0.255 ;
      RECT 0.836 0.225 0.866 0.255 ;
      RECT 0.614 0.225 0.644 0.255 ;
      RECT 0.466 0.225 0.496 0.255 ;
      RECT 2.02 0.165 2.05 0.195 ;
      RECT 1.65 0.165 1.68 0.195 ;
      RECT 0.91 0.105 0.94 0.135 ;
      RECT 0.54 0.105 0.57 0.135 ;
    LAYER NWELL ;
      RECT -0.074 0.3 2.294 0.6 ;
    LAYER DIFF ;
      RECT 0.518 0.45 2.146 0.55 ;
      RECT 0.074 0.45 0.444 0.55 ;
      RECT 0.074 0.05 2.146 0.15 ;
    LAYER PO ;
      RECT 2.213 0 2.227 0.6 ;
      RECT 2.139 0 2.153 0.6 ;
      RECT 2.065 0 2.079 0.6 ;
      RECT 1.991 0 2.005 0.6 ;
      RECT 1.917 0 1.931 0.6 ;
      RECT 1.843 0 1.857 0.6 ;
      RECT 1.769 0 1.783 0.6 ;
      RECT 1.695 0 1.709 0.6 ;
      RECT 1.621 0 1.635 0.6 ;
      RECT 1.547 0 1.561 0.6 ;
      RECT 1.473 0 1.487 0.6 ;
      RECT 1.399 0 1.413 0.6 ;
      RECT 1.325 0 1.339 0.6 ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_FSDPSYNSBQ_V2LP_0P5

MACRO SAEDRVT14_FDP_V2LP_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.554 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.15 0.128 0.446 ;
        RECT MASK 1 0.094 0.15 0.128 0.446 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.28 0.285 1.31 0.315 ;
      LAYER M2 ;
        RECT 1.038 0.283 1.401 0.317 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.058 0.405 1.088 0.435 ;
      LAYER M2 ;
        RECT 0.961 0.403 1.185 0.437 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.426 0.091 1.46 0.507 ;
        RECT MASK 1 1.426 0.091 1.46 0.507 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.596 0.647 ;
        RECT MASK 1 -0.042 0.553 1.596 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.046 1.596 0.048 ;
        RECT MASK 1 -0.042 -0.046 1.596 0.048 ;
    END
  END VSS
  OBS
    LAYER M2 ;
      RECT MASK 1 0.16 0.343 1.26 0.377 ;
      RECT MASK 1 0.294 0.223 1.192 0.257 ;
    LAYER VIA1 ;
      RECT 1.206 0.345 1.236 0.375 ;
      RECT 0.614 0.345 0.644 0.375 ;
      RECT 0.17 0.345 0.2 0.375 ;
      RECT 0.91 0.285 0.94 0.315 ;
      RECT 0.762 0.285 0.792 0.315 ;
      RECT 0.497 0.285 0.527 0.315 ;
      RECT 0.244 0.285 0.274 0.315 ;
      RECT 1.132 0.225 1.162 0.255 ;
      RECT 0.688 0.225 0.718 0.255 ;
      RECT 0.318 0.225 0.348 0.255 ;
      RECT 1.354 0.165 1.384 0.195 ;
      RECT 0.836 0.165 0.866 0.195 ;
    LAYER M1 ;
      RECT MASK 1 1.056 0.091 1.09 0.507 ;
      RECT MASK 1 0.316 0.41 0.35 0.507 ;
      RECT MASK 1 0.242 0.376 0.35 0.41 ;
      RECT MASK 1 0.242 0.091 0.276 0.376 ;
      RECT MASK 1 1.204 0.464 1.335 0.498 ;
      RECT MASK 1 1.204 0.137 1.238 0.464 ;
      RECT MASK 1 1.204 0.103 1.335 0.137 ;
      RECT MASK 1 0.67 0.464 0.868 0.498 ;
      RECT MASK 1 0.834 0.138 0.868 0.464 ;
      RECT MASK 1 0.59 0.104 0.868 0.138 ;
      RECT MASK 1 0.419 0.464 0.594 0.498 ;
      RECT MASK 1 0.419 0.222 0.453 0.464 ;
      RECT MASK 1 0.419 0.188 0.572 0.222 ;
      RECT MASK 1 1.13 0.123 1.164 0.477 ;
      RECT MASK 1 0.908 0.315 0.942 0.477 ;
      RECT MASK 1 0.908 0.281 1.013 0.315 ;
      RECT MASK 1 0.908 0.123 0.942 0.281 ;
      RECT MASK 1 0.168 0.233 0.202 0.477 ;
      RECT MASK 1 1.352 0.163 1.386 0.424 ;
      RECT MASK 1 1.278 0.256 1.312 0.424 ;
      RECT MASK 1 0.495 0.263 0.529 0.424 ;
      RECT MASK 1 0.612 0.206 0.646 0.422 ;
      RECT MASK 1 0.76 0.206 0.794 0.392 ;
      RECT MASK 1 0.686 0.206 0.72 0.392 ;
      RECT MASK 1 0.316 0.165 0.35 0.326 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.628 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 1.48 0.55 ;
      RECT 0.962 0.35 1.11 0.45 ;
      RECT 1.332 0.35 1.48 0.45 ;
      RECT 0.962 0.15 1.11 0.25 ;
      RECT 1.332 0.15 1.48 0.25 ;
      RECT 0.074 0.05 1.48 0.15 ;
    LAYER PO ;
      RECT 1.547 0 1.561 0.6 ;
      RECT 1.473 0 1.487 0.6 ;
      RECT 1.399 0 1.413 0.6 ;
      RECT 1.325 0 1.339 0.6 ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_FDP_V2LP_1

MACRO SAEDRVT14_FDPCBQ_V2LP_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.628 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.163 0.276 0.424 ;
        RECT 0.242 0.163 0.276 0.424 ;
    END
  END D
  PIN RS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.109 0.225 0.139 0.255 ;
      LAYER M2 ;
        RECT -0.028 0.223 0.164 0.257 ;
        RECT MASK 1 -0.028 0.223 0.164 0.257 ;
    END
  END RS
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.354 0.165 1.384 0.195 ;
      LAYER M2 ;
        RECT 1.034 0.163 1.386 0.197 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 1.5 0.093 1.534 0.507 ;
        RECT 1.5 0.093 1.534 0.507 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.67 0.647 ;
        RECT MASK 1 -0.042 0.553 1.67 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 -0.047 1.67 0.047 ;
        RECT -0.042 -0.047 1.67 0.047 ;
    END
  END VSS
  OBS
    LAYER M2 ;
      RECT MASK 1 0.506 0.343 1.266 0.377 ;
      RECT MASK 1 0.368 0.223 1.312 0.257 ;
    LAYER VIA1 ;
      RECT 1.206 0.345 1.236 0.375 ;
      RECT 0.803 0.345 0.833 0.375 ;
      RECT 0.54 0.345 0.57 0.375 ;
      RECT 1.428 0.285 1.458 0.315 ;
      RECT 1.132 0.285 1.162 0.315 ;
      RECT 0.984 0.285 1.014 0.315 ;
      RECT 0.701 0.285 0.731 0.315 ;
      RECT 0.466 0.285 0.496 0.315 ;
      RECT 1.28 0.225 1.31 0.255 ;
      RECT 0.883 0.225 0.913 0.255 ;
      RECT 0.392 0.225 0.422 0.255 ;
    LAYER M1 ;
      RECT MASK 1 1.278 0.464 1.386 0.498 ;
      RECT MASK 1 1.278 0.136 1.312 0.464 ;
      RECT MASK 1 1.278 0.102 1.407 0.136 ;
      RECT MASK 1 0.891 0.464 1.09 0.498 ;
      RECT MASK 1 1.056 0.136 1.09 0.464 ;
      RECT MASK 1 0.811 0.102 1.09 0.136 ;
      RECT MASK 1 0.612 0.464 0.812 0.498 ;
      RECT MASK 1 0.612 0.21 0.646 0.464 ;
      RECT MASK 1 0.612 0.176 0.806 0.21 ;
      RECT MASK 1 0.39 0.411 0.424 0.498 ;
      RECT MASK 1 0.39 0.377 0.498 0.411 ;
      RECT MASK 1 0.464 0.102 0.498 0.377 ;
      RECT MASK 1 0.151 0.464 0.35 0.498 ;
      RECT MASK 1 0.311 0.392 0.35 0.464 ;
      RECT MASK 1 1.204 0.124 1.238 0.478 ;
      RECT MASK 1 0.538 0.233 0.572 0.477 ;
      RECT MASK 1 1.13 0.161 1.164 0.475 ;
      RECT MASK 1 1.426 0.205 1.46 0.434 ;
      RECT MASK 1 1.352 0.163 1.386 0.424 ;
      RECT MASK 1 0.801 0.263 0.835 0.424 ;
      RECT MASK 1 0.699 0.263 0.733 0.424 ;
      RECT MASK 1 0.982 0.176 1.016 0.392 ;
      RECT MASK 1 0.881 0.206 0.915 0.392 ;
      RECT MASK 1 0.107 0.163 0.141 0.326 ;
      RECT MASK 1 0.39 0.162 0.424 0.325 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.702 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 1.554 0.55 ;
      RECT 1.406 0.35 1.554 0.45 ;
      RECT 1.406 0.15 1.554 0.25 ;
      RECT 0.37 0.05 1.554 0.15 ;
      RECT 0.074 0.05 0.296 0.15 ;
    LAYER PO ;
      RECT 1.621 0 1.635 0.6 ;
      RECT 1.547 0 1.561 0.6 ;
      RECT 1.473 0 1.487 0.6 ;
      RECT 1.399 0 1.413 0.6 ;
      RECT 1.325 0 1.339 0.6 ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_FDPCBQ_V2LP_1

MACRO SAEDRVT14_FSDPQ_V2LP_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.85 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.464 0.194 0.498 0.418 ;
        RECT 0.464 0.194 0.498 0.418 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.118 0.202 0.313 ;
        RECT 0.168 0.118 0.202 0.313 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.196 0.424 0.418 ;
        RECT 0.39 0.196 0.424 0.418 ;
    END
  END SE
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.576 0.345 1.606 0.375 ;
      LAYER M2 ;
        RECT MASK 1 1.554 0.343 1.79 0.377 ;
        RECT 1.554 0.343 1.79 0.377 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 1.722 0.088 1.756 0.488 ;
        RECT 1.722 0.088 1.756 0.488 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.892 0.647 ;
        RECT MASK 1 -0.042 0.553 1.892 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.892 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.892 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.269 0.458 0.578 0.496 ;
      RECT MASK 1 0.544 0.139 0.578 0.458 ;
      RECT MASK 1 0.347 0.105 0.578 0.139 ;
      RECT MASK 1 1.427 0.118 1.461 0.458 ;
      RECT MASK 1 1.352 0.118 1.386 0.458 ;
      RECT MASK 1 0.618 0.224 0.652 0.458 ;
      RECT MASK 1 1.071 0.199 1.105 0.437 ;
      RECT MASK 1 0.953 0.263 0.999 0.42 ;
      RECT MASK 1 1.651 0.197 1.685 0.418 ;
      RECT MASK 1 1.589 0.163 1.685 0.197 ;
      RECT MASK 1 1.567 0.278 1.611 0.413 ;
      RECT MASK 1 1.213 0.199 1.247 0.377 ;
      RECT MASK 1 0.756 0.158 0.802 0.317 ;
    LAYER M2 ;
      RECT MASK 1 1.172 0.343 1.474 0.377 ;
      RECT MASK 1 0.686 0.343 1.051 0.377 ;
    LAYER VIA1 ;
      RECT 1.502 0.405 1.532 0.435 ;
      RECT 1.073 0.405 1.103 0.435 ;
      RECT 0.62 0.405 0.65 0.435 ;
      RECT 1.354 0.345 1.384 0.375 ;
      RECT 1.215 0.345 1.245 0.375 ;
      RECT 0.96 0.345 0.99 0.375 ;
      RECT 0.688 0.345 0.718 0.375 ;
      RECT 1.429 0.285 1.459 0.315 ;
      RECT 1.144 0.285 1.174 0.315 ;
      RECT 0.763 0.285 0.793 0.315 ;
      RECT 1.593 0.165 1.623 0.195 ;
      RECT 1.282 0.165 1.312 0.195 ;
    LAYER NWELL ;
      RECT -0.074 0.289 1.924 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 1.776 0.55 ;
      RECT 0.074 0.05 1.776 0.15 ;
    LAYER PO ;
      RECT 1.843 0 1.857 0.6 ;
      RECT 1.769 0 1.783 0.6 ;
      RECT 1.695 0 1.709 0.6 ;
      RECT 1.621 0 1.635 0.6 ;
      RECT 1.547 0 1.561 0.6 ;
      RECT 1.473 0 1.487 0.6 ;
      RECT 1.399 0 1.413 0.6 ;
      RECT 1.325 0 1.339 0.6 ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_FSDPQ_V2LP_0P5

MACRO SAEDRVT14_FDPQB_V2LP_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.406 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.112 0.128 0.488 ;
        RECT MASK 1 0.094 0.112 0.128 0.488 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.129 0.285 1.159 0.315 ;
      LAYER M2 ;
        RECT 1.086 0.283 1.323 0.317 ;
    END
  END CK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.3 0.405 1.33 0.435 ;
      LAYER M2 ;
        RECT 1.029 0.403 1.413 0.437 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.448 0.647 ;
        RECT MASK 1 -0.042 0.553 1.448 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.448 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.448 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 1.298 0.112 1.332 0.488 ;
      RECT MASK 1 1.059 0.45 1.198 0.488 ;
      RECT MASK 1 1.059 0.15 1.093 0.45 ;
      RECT MASK 1 1.059 0.112 1.196 0.15 ;
      RECT MASK 1 0.394 0.45 0.581 0.488 ;
      RECT MASK 1 0.394 0.215 0.44 0.45 ;
      RECT MASK 1 0.394 0.181 0.575 0.215 ;
      RECT MASK 1 0.24 0.454 0.34 0.488 ;
      RECT MASK 1 0.24 0.112 0.274 0.454 ;
      RECT MASK 1 0.916 0.118 0.95 0.458 ;
      RECT MASK 1 0.622 0.19 0.656 0.418 ;
      RECT MASK 1 0.768 0.199 0.802 0.377 ;
    LAYER M2 ;
      RECT MASK 1 0.164 0.343 1.168 0.377 ;
      RECT MASK 1 0.307 0.223 1.096 0.257 ;
    LAYER VIA1 ;
      RECT 1.061 0.345 1.091 0.375 ;
      RECT 0.624 0.345 0.654 0.375 ;
      RECT 0.172 0.345 0.202 0.375 ;
      RECT 0.918 0.285 0.948 0.315 ;
      RECT 0.77 0.285 0.8 0.315 ;
      RECT 0.495 0.285 0.525 0.315 ;
      RECT 0.242 0.285 0.272 0.315 ;
      RECT 0.992 0.225 1.022 0.255 ;
      RECT 0.699 0.225 0.729 0.255 ;
      RECT 0.314 0.225 0.344 0.255 ;
      RECT 1.231 0.165 1.261 0.195 ;
      RECT 0.842 0.165 0.872 0.195 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.48 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 1.332 0.55 ;
      RECT 0.074 0.05 1.332 0.15 ;
    LAYER PO ;
      RECT 1.399 0 1.413 0.6 ;
      RECT 1.325 0 1.339 0.6 ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_FDPQB_V2LP_0P5

MACRO SAEDRVT14_FDPQB_V2LP_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.406 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.112 0.128 0.488 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.129 0.285 1.159 0.315 ;
      LAYER M2 ;
        RECT 1.086 0.283 1.323 0.317 ;
    END
  END CK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.3 0.405 1.33 0.435 ;
      LAYER M2 ;
        RECT 1.029 0.403 1.413 0.437 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.448 0.647 ;
        RECT MASK 1 -0.042 0.553 1.448 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.448 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.448 0.047 ;
    END
  END VSS
  OBS
    LAYER M2 ;
      RECT MASK 1 0.164 0.343 1.168 0.377 ;
      RECT MASK 1 0.306 0.223 1.096 0.257 ;
    LAYER VIA1 ;
      RECT 1.061 0.345 1.091 0.375 ;
      RECT 0.624 0.345 0.654 0.375 ;
      RECT 0.172 0.345 0.202 0.375 ;
      RECT 0.918 0.285 0.948 0.315 ;
      RECT 0.77 0.285 0.8 0.315 ;
      RECT 0.495 0.285 0.525 0.315 ;
      RECT 0.242 0.285 0.272 0.315 ;
      RECT 0.992 0.225 1.022 0.255 ;
      RECT 0.699 0.225 0.729 0.255 ;
      RECT 0.314 0.225 0.344 0.255 ;
      RECT 1.221 0.165 1.251 0.195 ;
      RECT 0.842 0.165 0.872 0.195 ;
    LAYER M1 ;
      RECT MASK 1 0.99 0.118 1.024 0.458 ;
      RECT MASK 1 0.916 0.118 0.95 0.458 ;
      RECT MASK 1 0.17 0.224 0.204 0.458 ;
      RECT MASK 1 1.219 0.163 1.253 0.423 ;
      RECT MASK 1 0.622 0.199 0.656 0.418 ;
      RECT MASK 1 1.127 0.25 1.161 0.416 ;
      RECT MASK 1 0.488 0.263 0.534 0.414 ;
      RECT MASK 1 0.307 0.158 0.353 0.409 ;
      RECT MASK 1 0.768 0.199 0.802 0.377 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.48 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 1.332 0.55 ;
      RECT 1.184 0.35 1.332 0.45 ;
      RECT 1.184 0.15 1.332 0.25 ;
      RECT 0.074 0.05 1.332 0.15 ;
    LAYER PO ;
      RECT 1.399 0 1.413 0.6 ;
      RECT 1.325 0 1.339 0.6 ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_FDPQB_V2LP_1

MACRO SAEDRVT14_FSDPSYNRBQ_V2LP_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.072 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN RD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.171 0.128 0.365 ;
        RECT 0.094 0.171 0.128 0.365 ;
    END
  END RD
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.176 0.276 0.418 ;
        RECT MASK 1 0.242 0.176 0.276 0.418 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.614 0.345 0.644 0.375 ;
      LAYER M2 ;
        RECT 0.409 0.343 0.691 0.377 ;
        RECT MASK 1 0.409 0.343 0.691 0.377 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.54 0.225 0.57 0.255 ;
      LAYER M2 ;
        RECT 0.409 0.223 0.691 0.257 ;
        RECT MASK 1 0.409 0.223 0.691 0.257 ;
    END
  END SE
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.657 0.285 1.687 0.315 ;
      LAYER M2 ;
        RECT 1.654 0.283 1.95 0.317 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.944 0.088 1.978 0.504 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 2.114 0.647 ;
        RECT MASK 1 -0.042 0.553 2.114 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 -0.047 2.114 0.047 ;
        RECT -0.042 -0.047 2.114 0.047 ;
    END
  END VSS
  OBS
    LAYER M2 ;
      RECT MASK 1 0.932 0.223 1.846 0.257 ;
      RECT MASK 1 0.329 0.103 0.818 0.137 ;
    LAYER VIA1 ;
      RECT 1.724 0.405 1.754 0.435 ;
      RECT 1.28 0.405 1.31 0.435 ;
      RECT 0.836 0.405 0.866 0.435 ;
      RECT 1.576 0.285 1.606 0.315 ;
      RECT 1.428 0.285 1.458 0.315 ;
      RECT 1.148 0.285 1.178 0.315 ;
      RECT 0.91 0.285 0.94 0.315 ;
      RECT 1.798 0.225 1.828 0.255 ;
      RECT 1.354 0.225 1.384 0.255 ;
      RECT 0.984 0.225 1.014 0.255 ;
      RECT 1.872 0.165 1.902 0.195 ;
      RECT 1.502 0.165 1.532 0.195 ;
      RECT 0.688 0.165 0.718 0.195 ;
      RECT 0.466 0.165 0.496 0.195 ;
      RECT 0.318 0.165 0.348 0.195 ;
      RECT 0.762 0.105 0.792 0.135 ;
      RECT 0.392 0.105 0.422 0.135 ;
    LAYER M1 ;
      RECT MASK 1 1.574 0.118 1.608 0.458 ;
      RECT MASK 1 0.834 0.224 0.868 0.458 ;
      RECT MASK 1 0.612 0.263 0.646 0.458 ;
      RECT MASK 1 1.278 0.206 1.312 0.437 ;
      RECT MASK 1 1.655 0.219 1.689 0.422 ;
      RECT MASK 1 1.14 0.263 1.186 0.418 ;
      RECT MASK 1 1.87 0.163 1.904 0.409 ;
      RECT MASK 1 1.426 0.199 1.46 0.377 ;
      RECT MASK 1 0.316 0.163 0.35 0.357 ;
      RECT MASK 1 0.982 0.158 1.016 0.313 ;
      RECT MASK 1 0.464 0.118 0.498 0.313 ;
    LAYER NWELL ;
      RECT -0.074 0.3 2.146 0.6 ;
    LAYER DIFF ;
      RECT 0.37 0.45 1.998 0.55 ;
      RECT 0.074 0.45 0.296 0.55 ;
      RECT 0.074 0.05 1.998 0.15 ;
    LAYER PO ;
      RECT 2.065 0 2.079 0.6 ;
      RECT 1.991 0 2.005 0.6 ;
      RECT 1.917 0 1.931 0.6 ;
      RECT 1.843 0 1.857 0.6 ;
      RECT 1.769 0 1.783 0.6 ;
      RECT 1.695 0 1.709 0.6 ;
      RECT 1.621 0 1.635 0.6 ;
      RECT 1.547 0 1.561 0.6 ;
      RECT 1.473 0 1.487 0.6 ;
      RECT 1.399 0 1.413 0.6 ;
      RECT 1.325 0 1.339 0.6 ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_FSDPSYNRBQ_V2LP_0P5

MACRO SAEDRVT14_ND2B_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.518 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.267 0.128 0.415 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.163 0.424 0.437 ;
        RECT 0.39 0.163 0.424 0.437 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.102 0.35 0.507 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.56 0.647 ;
        RECT MASK 1 -0.042 0.553 0.56 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.56 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.56 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.144 0.443 0.276 0.477 ;
      RECT MASK 1 0.242 0.21 0.276 0.443 ;
      RECT MASK 1 0.142 0.176 0.276 0.21 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.592 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.444 0.55 ;
      RECT 0.074 0.05 0.444 0.15 ;
    LAYER PO ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_ND2B_U_0P5

MACRO SAEDRVT14_AO221_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.814 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.207 0.285 0.237 0.315 ;
      LAYER M2 ;
        RECT 0.085 0.283 0.321 0.317 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.089 0.128 0.289 ;
        RECT 0.094 0.089 0.128 0.289 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.316 0.168 0.35 0.357 ;
        RECT 0.316 0.168 0.35 0.357 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.168 0.424 0.357 ;
        RECT 0.39 0.168 0.424 0.357 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.526 0.225 0.556 0.255 ;
      LAYER M2 ;
        RECT 0.491 0.223 0.679 0.257 ;
        RECT MASK 1 0.491 0.223 0.679 0.257 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.686 0.119 0.72 0.459 ;
        RECT MASK 1 0.686 0.119 0.72 0.459 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.856 0.647 ;
        RECT MASK 1 -0.042 0.553 0.856 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.856 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.856 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.54 0.459 0.643 0.497 ;
      RECT MASK 1 0.609 0.142 0.643 0.459 ;
      RECT MASK 1 0.228 0.104 0.643 0.142 ;
      RECT MASK 1 0.103 0.459 0.46 0.497 ;
      RECT MASK 1 0.103 0.37 0.141 0.459 ;
      RECT MASK 1 0.304 0.383 0.544 0.417 ;
      RECT MASK 1 0.205 0.182 0.239 0.384 ;
      RECT MASK 1 0.519 0.204 0.565 0.343 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.888 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.74 0.55 ;
      RECT 0.074 0.4 0.592 0.45 ;
      RECT 0.074 0.05 0.74 0.15 ;
    LAYER PO ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AO221_0P5

MACRO SAEDRVT14_INV_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.296 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.159 0.128 0.419 ;
        RECT 0.094 0.159 0.128 0.419 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.089 0.202 0.489 ;
        RECT 0.168 0.089 0.202 0.489 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 0.553 0.338 0.647 ;
        RECT -0.042 0.553 0.338 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 -0.048 0.338 0.046 ;
        RECT -0.042 -0.048 0.338 0.046 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.3 0.37 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.35 0.222 0.55 ;
      RECT 0.074 0.05 0.222 0.25 ;
    LAYER PO ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_INV_1

MACRO SAEDRVT14_ND2_CDC_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.37 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.165 0.128 0.435 ;
        RECT MASK 1 0.094 0.165 0.128 0.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.274 0.276 0.477 ;
        RECT 0.242 0.274 0.276 0.477 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.224 0.202 0.509 ;
        RECT MASK 1 0.168 0.188 0.276 0.224 ;
        RECT MASK 1 0.242 0.091 0.276 0.188 ;
        RECT 0.168 0.188 0.202 0.509 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.55 0.412 0.647 ;
        RECT MASK 1 -0.042 0.55 0.412 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.412 0.05 ;
        RECT MASK 1 -0.042 -0.047 0.412 0.05 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.3 0.444 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.296 0.55 ;
      RECT 0.074 0.05 0.296 0.25 ;
    LAYER PO ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_ND2_CDC_0P5

MACRO SAEDRVT14_OR3_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.592 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.316 0.216 0.35 0.418 ;
        RECT 0.316 0.216 0.35 0.418 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.216 0.276 0.418 ;
        RECT 0.242 0.216 0.276 0.418 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.199 0.128 0.488 ;
        RECT 0.094 0.199 0.128 0.488 ;
    END
  END A3
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.464 0.118 0.498 0.458 ;
        RECT 0.464 0.118 0.498 0.458 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.634 0.647 ;
        RECT MASK 1 -0.042 0.553 0.634 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.634 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.634 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.304 0.458 0.424 0.496 ;
      RECT MASK 1 0.39 0.136 0.424 0.458 ;
      RECT MASK 1 0.15 0.102 0.424 0.136 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.666 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.518 0.55 ;
      RECT 0.155 0.4 0.369 0.45 ;
      RECT 0.074 0.05 0.518 0.15 ;
    LAYER PO ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OR3_0P5

MACRO SAEDRVT14_INV_0P75
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.296 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.159 0.128 0.419 ;
        RECT MASK 1 0.094 0.159 0.128 0.419 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.089 0.202 0.489 ;
        RECT MASK 1 0.168 0.089 0.202 0.489 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.338 0.647 ;
        RECT MASK 1 -0.042 0.553 0.338 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.048 0.338 0.046 ;
        RECT MASK 1 -0.042 -0.048 0.338 0.046 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.3 0.37 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.35 0.222 0.5 ;
      RECT 0.074 0.05 0.222 0.2 ;
    LAYER PO ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_INV_0P75

MACRO SAEDRVT14_INV_S_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.296 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.159 0.128 0.419 ;
        RECT 0.094 0.159 0.128 0.419 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.089 0.202 0.489 ;
        RECT 0.168 0.089 0.202 0.489 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.338 0.647 ;
        RECT MASK 1 -0.042 0.553 0.338 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.048 0.338 0.046 ;
        RECT MASK 1 -0.042 -0.048 0.338 0.046 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.078 0.3 0.37 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.222 0.5 ;
      RECT 0.074 0.05 0.222 0.15 ;
    LAYER PO ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_INV_S_0P5

MACRO SAEDRVT14_OA21B_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.592 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.199 0.276 0.386 ;
        RECT MASK 1 0.242 0.199 0.276 0.386 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.115 0.225 0.145 0.255 ;
      LAYER M2 ;
        RECT MASK 1 -0.035 0.223 0.147 0.257 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.475 0.105 0.505 0.135 ;
      LAYER M2 ;
        RECT MASK 1 0.473 0.103 0.622 0.137 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.401 0.165 0.431 0.195 ;
      LAYER M2 ;
        RECT 0.26 0.163 0.434 0.197 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 0.553 0.634 0.647 ;
        RECT -0.042 0.553 0.634 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.634 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.634 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.459 0.395 0.499 0.488 ;
      RECT MASK 1 0.399 0.361 0.499 0.395 ;
      RECT MASK 1 0.399 0.088 0.433 0.361 ;
      RECT MASK 1 0.216 0.422 0.359 0.46 ;
      RECT MASK 1 0.325 0.154 0.359 0.422 ;
      RECT MASK 1 0.138 0.112 0.359 0.154 ;
      RECT MASK 1 0.112 0.199 0.147 0.442 ;
      RECT MASK 1 0.473 0.103 0.507 0.313 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.666 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.35 0.518 0.55 ;
      RECT 0.074 0.05 0.518 0.15 ;
    LAYER PO ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OA21B_1

MACRO SAEDRVT14_OAI22_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.518 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.199 0.276 0.377 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.392 0.285 0.422 0.315 ;
      LAYER M2 ;
        RECT 0.276 0.283 0.43 0.317 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.158 0.202 0.354 ;
        RECT MASK 1 0.168 0.158 0.202 0.354 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.263 0.128 0.488 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.158 0.35 0.46 ;
        RECT MASK 1 0.225 0.422 0.35 0.46 ;
        RECT MASK 1 0.316 0.158 0.35 0.422 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.56 0.647 ;
        RECT MASK 1 -0.042 0.553 0.56 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.56 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.56 0.047 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.3 0.592 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.464 0.55 ;
      RECT 0.074 0.05 0.464 0.15 ;
    LAYER PO ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OAI22_0P5

MACRO SAEDRVT14_AOI21_0P75
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.444 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.222 0.202 0.414 ;
        RECT 0.168 0.222 0.202 0.414 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.199 0.128 0.377 ;
        RECT 0.094 0.199 0.128 0.377 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.199 0.276 0.377 ;
        RECT 0.242 0.199 0.276 0.377 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.316 0.146 0.35 0.415 ;
        RECT MASK 1 0.23 0.112 0.35 0.146 ;
        RECT 0.316 0.112 0.35 0.415 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.486 0.647 ;
        RECT MASK 1 -0.042 0.553 0.486 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.486 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.486 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.094 0.454 0.304 0.488 ;
      RECT MASK 1 0.094 0.417 0.128 0.454 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.518 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.37 0.55 ;
      RECT 0.074 0.35 0.215 0.4 ;
      RECT 0.155 0.2 0.289 0.25 ;
      RECT 0.074 0.15 0.289 0.2 ;
      RECT 0.074 0.05 0.37 0.15 ;
    LAYER PO ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AOI21_0P75

MACRO SAEDRVT14_AO32_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.74 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.245 0.345 0.275 0.375 ;
      LAYER M2 ;
        RECT MASK 1 0.057 0.343 0.277 0.377 ;
        RECT 0.057 0.343 0.277 0.377 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.102 0.202 0.377 ;
        RECT MASK 1 0.168 0.102 0.202 0.377 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.121 0.128 0.381 ;
        RECT 0.094 0.121 0.128 0.381 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.324 0.285 0.354 0.315 ;
      LAYER M2 ;
        RECT 0.268 0.283 0.43 0.317 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.456 0.225 0.486 0.255 ;
      LAYER M2 ;
        RECT MASK 1 0.4 0.223 0.562 0.257 ;
        RECT 0.4 0.223 0.562 0.257 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.614 0.105 0.644 0.135 ;
      LAYER M2 ;
        RECT 0.555 0.103 0.834 0.137 ;
        RECT MASK 1 0.555 0.103 0.834 0.137 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.782 0.647 ;
        RECT MASK 1 -0.042 0.553 0.782 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.782 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.782 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.15 0.46 0.544 0.498 ;
      RECT MASK 1 0.612 0.088 0.646 0.488 ;
      RECT MASK 1 0.358 0.386 0.572 0.42 ;
      RECT MASK 1 0.538 0.148 0.572 0.386 ;
      RECT MASK 1 0.28 0.11 0.572 0.148 ;
      RECT MASK 1 0.243 0.224 0.277 0.418 ;
      RECT MASK 1 0.451 0.193 0.497 0.346 ;
      RECT MASK 1 0.317 0.193 0.363 0.346 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.814 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.666 0.55 ;
      RECT 0.229 0.2 0.303 0.25 ;
      RECT 0.155 0.15 0.377 0.2 ;
      RECT 0.074 0.05 0.666 0.15 ;
    LAYER PO ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
      RECT 0.733 0 0.747 0.59 ;
  END
END SAEDRVT14_AO32_U_0P5

MACRO SAEDRVT14_OR3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.592 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.316 0.216 0.35 0.418 ;
        RECT 0.316 0.216 0.35 0.418 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.216 0.276 0.418 ;
        RECT 0.242 0.216 0.276 0.418 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.199 0.128 0.488 ;
        RECT 0.094 0.199 0.128 0.488 ;
    END
  END A3
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.464 0.118 0.498 0.458 ;
        RECT 0.464 0.118 0.498 0.458 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.634 0.647 ;
        RECT MASK 1 -0.042 0.553 0.634 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.634 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.634 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.304 0.458 0.424 0.496 ;
      RECT MASK 1 0.39 0.136 0.424 0.458 ;
      RECT MASK 1 0.15 0.102 0.424 0.136 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.666 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.518 0.55 ;
      RECT 0.369 0.35 0.518 0.4 ;
      RECT 0.37 0.15 0.518 0.25 ;
      RECT 0.074 0.05 0.518 0.15 ;
    LAYER PO ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OR3_1

MACRO SAEDRVT14_INV_PS_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.296 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.106 0.128 0.317 ;
        RECT 0.094 0.106 0.128 0.317 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.118 0.202 0.378 ;
        RECT 0.168 0.118 0.202 0.378 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.597 0.338 0.691 ;
        RECT MASK 1 -0.042 0.597 0.338 0.691 ;
    END
  END VDD
  PIN VDDR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.096 0.463 0.126 0.493 ;
      LAYER M2 ;
        RECT 0.094 0.457 0.2 0.543 ;
        RECT MASK 1 0.094 0.457 0.2 0.543 ;
    END
  END VDDR
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 -0.047 0.338 0.047 ;
        RECT -0.042 -0.047 0.338 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.094 0.464 0.2 0.498 ;
      RECT MASK 1 0.094 0.357 0.128 0.464 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.37 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.35 0.222 0.55 ;
      RECT 0.074 0.05 0.222 0.25 ;
    LAYER PO ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_INV_PS_1

MACRO SAEDRVT14_NR2_MM_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.37 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.123 0.276 0.349 ;
        RECT 0.242 0.123 0.276 0.349 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.165 0.128 0.435 ;
        RECT 0.094 0.165 0.128 0.435 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.091 0.202 0.441 ;
        RECT MASK 1 0.24 0.441 0.274 0.509 ;
        RECT MASK 1 0.168 0.404 0.274 0.441 ;
        RECT MASK 1 0.168 0.091 0.202 0.404 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.55 0.412 0.647 ;
        RECT MASK 1 -0.042 0.55 0.412 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.412 0.05 ;
        RECT MASK 1 -0.042 -0.047 0.412 0.05 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.299 0.444 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.35 0.308 0.55 ;
      RECT 0.074 0.05 0.308 0.2 ;
    LAYER PO ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_NR2_MM_1

MACRO SAEDRVT14_AN2_MM_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.518 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.186 0.202 0.412 ;
        RECT 0.168 0.186 0.202 0.412 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.096 0.225 0.126 0.255 ;
      LAYER M2 ;
        RECT 0.029 0.223 0.219 0.257 ;
        RECT MASK 1 0.029 0.223 0.219 0.257 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.123 0.424 0.477 ;
        RECT 0.39 0.123 0.424 0.477 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.56 0.647 ;
        RECT MASK 1 -0.042 0.553 0.56 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.56 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.56 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.094 0.091 0.128 0.334 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.592 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.444 0.55 ;
      RECT 0.296 0.35 0.444 0.45 ;
      RECT 0.296 0.2 0.444 0.25 ;
      RECT 0.074 0.05 0.444 0.2 ;
    LAYER PO ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AN2_MM_1

MACRO SAEDRVT14_INV_S_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.296 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.159 0.128 0.419 ;
        RECT 0.094 0.159 0.128 0.419 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.089 0.202 0.489 ;
        RECT 0.168 0.089 0.202 0.489 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.338 0.647 ;
        RECT MASK 1 -0.042 0.553 0.338 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 -0.048 0.338 0.046 ;
        RECT -0.042 -0.048 0.338 0.046 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.078 0.3 0.37 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.35 0.222 0.55 ;
      RECT 0.074 0.05 0.222 0.25 ;
    LAYER PO ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_INV_S_1

MACRO SAEDRVT14_NR3_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.74 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.199 0.276 0.442 ;
        RECT MASK 1 0.242 0.199 0.276 0.442 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.199 0.202 0.502 ;
        RECT MASK 1 0.168 0.199 0.202 0.502 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.2 0.128 0.441 ;
        RECT MASK 1 0.094 0.2 0.128 0.441 ;
    END
  END A3
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.099 0.646 0.503 ;
        RECT MASK 1 0.612 0.099 0.646 0.503 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.782 0.647 ;
        RECT MASK 1 -0.042 0.553 0.782 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 -0.047 0.782 0.047 ;
        RECT -0.042 -0.047 0.782 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.437 0.454 0.572 0.488 ;
      RECT MASK 1 0.538 0.146 0.572 0.454 ;
      RECT MASK 1 0.437 0.112 0.572 0.146 ;
      RECT MASK 1 0.316 0.316 0.35 0.488 ;
      RECT MASK 1 0.427 0.316 0.461 0.414 ;
      RECT MASK 1 0.316 0.282 0.461 0.316 ;
      RECT MASK 1 0.427 0.186 0.461 0.282 ;
      RECT MASK 1 0.316 0.146 0.35 0.282 ;
      RECT MASK 1 0.146 0.112 0.35 0.146 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.814 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.666 0.55 ;
      RECT 0.074 0.35 0.37 0.45 ;
      RECT 0.518 0.35 0.666 0.45 ;
      RECT 0.074 0.2 0.289 0.25 ;
      RECT 0.518 0.2 0.666 0.25 ;
      RECT 0.074 0.05 0.666 0.2 ;
    LAYER PO ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_NR3_1

MACRO SAEDRVT14_OA31_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.666 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.185 0.276 0.352 ;
        RECT 0.242 0.185 0.276 0.352 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.199 0.202 0.488 ;
        RECT 0.168 0.199 0.202 0.488 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.185 0.128 0.418 ;
        RECT 0.094 0.185 0.128 0.418 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.24 0.424 0.396 ;
        RECT 0.39 0.24 0.424 0.396 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.538 0.088 0.572 0.488 ;
        RECT 0.538 0.088 0.572 0.488 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.708 0.647 ;
        RECT MASK 1 -0.042 0.553 0.708 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.708 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.708 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.306 0.422 0.512 0.46 ;
      RECT MASK 1 0.478 0.214 0.512 0.422 ;
      RECT MASK 1 0.382 0.18 0.512 0.214 ;
      RECT MASK 1 0.15 0.102 0.388 0.14 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.74 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.592 0.55 ;
      RECT 0.444 0.35 0.592 0.4 ;
      RECT 0.444 0.2 0.592 0.25 ;
      RECT 0.074 0.05 0.592 0.2 ;
    LAYER PO ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OA31_1

MACRO SAEDRVT14_AN3_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.592 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.291 0.345 0.321 0.375 ;
      LAYER M2 ;
        RECT 0.281 0.343 0.458 0.377 ;
        RECT MASK 1 0.281 0.343 0.458 0.377 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.215 0.225 0.245 0.255 ;
      LAYER M2 ;
        RECT MASK 1 0.191 0.223 0.346 0.257 ;
        RECT 0.212 0.223 0.323 0.257 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.115 0.165 0.145 0.195 ;
      LAYER M2 ;
        RECT 0.03 0.163 0.165 0.197 ;
    END
  END A3
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.464 0.119 0.498 0.459 ;
        RECT MASK 1 0.464 0.119 0.498 0.459 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.634 0.647 ;
        RECT MASK 1 -0.042 0.553 0.634 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.634 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.634 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.15 0.45 0.424 0.488 ;
      RECT MASK 1 0.39 0.148 0.424 0.45 ;
      RECT MASK 1 0.304 0.114 0.424 0.148 ;
      RECT MASK 1 0.289 0.202 0.323 0.41 ;
      RECT MASK 1 0.213 0.159 0.247 0.409 ;
      RECT MASK 1 0.113 0.112 0.147 0.378 ;
    LAYER NWELL ;
      RECT -0.074 0.289 0.666 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.518 0.55 ;
      RECT 0.37 0.4 0.518 0.45 ;
      RECT 0.289 0.15 0.37 0.2 ;
      RECT 0.074 0.05 0.518 0.15 ;
    LAYER PO ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AN3_0P5

MACRO SAEDRVT14_OR4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.666 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.37 0.225 0.4 0.255 ;
      LAYER M2 ;
        RECT MASK 1 0.356 0.223 0.599 0.257 ;
        RECT 0.356 0.223 0.599 0.257 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.27 0.285 0.3 0.315 ;
      LAYER M2 ;
        RECT 0.262 0.283 0.461 0.317 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.192 0.345 0.222 0.375 ;
      LAYER M2 ;
        RECT 0.155 0.343 0.334 0.377 ;
        RECT MASK 1 0.155 0.343 0.334 0.377 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.114 0.405 0.144 0.435 ;
      LAYER M2 ;
        RECT 0.007 0.403 0.162 0.437 ;
    END
  END A4
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.538 0.118 0.572 0.458 ;
        RECT MASK 1 0.538 0.118 0.572 0.458 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.708 0.647 ;
        RECT MASK 1 -0.042 0.553 0.708 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.708 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.708 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.382 0.458 0.498 0.496 ;
      RECT MASK 1 0.464 0.136 0.498 0.458 ;
      RECT MASK 1 0.15 0.102 0.498 0.136 ;
      RECT MASK 1 0.268 0.199 0.302 0.488 ;
      RECT MASK 1 0.112 0.199 0.146 0.488 ;
      RECT MASK 1 0.368 0.176 0.402 0.418 ;
      RECT MASK 1 0.19 0.176 0.224 0.418 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.74 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.592 0.55 ;
      RECT 0.289 0.35 0.592 0.4 ;
      RECT 0.444 0.15 0.592 0.25 ;
      RECT 0.074 0.05 0.592 0.15 ;
    LAYER PO ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OR4_1

MACRO SAEDRVT14_INV_S_0P75
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.296 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.159 0.128 0.419 ;
        RECT 0.094 0.159 0.128 0.419 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.089 0.202 0.489 ;
        RECT MASK 1 0.168 0.089 0.202 0.489 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 0.553 0.338 0.647 ;
        RECT -0.042 0.553 0.338 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 -0.048 0.338 0.046 ;
        RECT -0.042 -0.048 0.338 0.046 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.078 0.3 0.37 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.35 0.222 0.5 ;
      RECT 0.074 0.05 0.222 0.2 ;
    LAYER PO ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_INV_S_0P75

MACRO SAEDRVT14_AO21_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.592 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.19 0.202 0.402 ;
        RECT MASK 1 0.168 0.19 0.202 0.402 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.112 0.128 0.288 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.19 0.276 0.382 ;
        RECT MASK 1 0.242 0.19 0.276 0.382 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.464 0.118 0.498 0.458 ;
        RECT MASK 1 0.464 0.118 0.498 0.458 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.635 0.647 ;
        RECT MASK 1 -0.042 0.553 0.635 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.635 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.635 0.047 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.3 0.667 0.6 ;
    LAYER DIFF ;
      RECT 0.075 0.45 0.519 0.55 ;
      RECT 0.075 0.05 0.519 0.15 ;
    LAYER PO ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AO21_U_0P5

MACRO SAEDRVT14_AN4_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.666 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 0.19 0.424 0.41 ;
        RECT MASK 1 0.39 0.19 0.424 0.41 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.112 0.35 0.377 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.165 0.276 0.41 ;
        RECT MASK 1 0.242 0.165 0.276 0.41 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.112 0.128 0.377 ;
    END
  END A4
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.533 0.165 0.563 0.195 ;
      LAYER M2 ;
        RECT 0.499 0.163 0.653 0.197 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.708 0.647 ;
        RECT MASK 1 -0.042 0.553 0.708 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.708 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.708 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.531 0.118 0.565 0.458 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.74 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.596 0.55 ;
      RECT 0.444 0.4 0.596 0.45 ;
      RECT 0.229 0.15 0.444 0.2 ;
      RECT 0.074 0.05 0.592 0.15 ;
    LAYER PO ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AN4_0P5

MACRO SAEDRVT14_MUX2_MM_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.74 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.123 0.202 0.326 ;
        RECT 0.168 0.123 0.202 0.326 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.464 0.176 0.498 0.424 ;
        RECT MASK 1 0.464 0.176 0.498 0.424 ;
    END
  END D1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.176 0.424 0.424 ;
        RECT 0.39 0.176 0.424 0.424 ;
    END
  END S
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.123 0.646 0.477 ;
        RECT MASK 1 0.612 0.123 0.646 0.477 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.786 0.647 ;
        RECT MASK 1 -0.042 0.553 0.786 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.786 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.786 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.366 0.464 0.572 0.498 ;
      RECT MASK 1 0.538 0.136 0.572 0.464 ;
      RECT MASK 1 0.292 0.102 0.572 0.136 ;
      RECT MASK 1 0.094 0.41 0.128 0.498 ;
      RECT MASK 1 0.094 0.376 0.296 0.41 ;
      RECT MASK 1 0.094 0.102 0.128 0.376 ;
      RECT MASK 1 0.262 0.206 0.296 0.376 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.818 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.67 0.55 ;
      RECT 0.074 0.05 0.67 0.15 ;
    LAYER PO ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_MUX2_MM_0P5

MACRO SAEDRVT14_AO21B_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.592 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.228 0.276 0.378 ;
        RECT MASK 1 0.242 0.228 0.276 0.378 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.089 0.128 0.378 ;
        RECT MASK 1 0.094 0.089 0.128 0.378 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.464 0.264 0.498 0.459 ;
        RECT 0.464 0.264 0.498 0.459 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.216 0.424 0.489 ;
        RECT MASK 1 0.39 0.182 0.499 0.216 ;
        RECT MASK 1 0.461 0.089 0.499 0.182 ;
        RECT 0.39 0.182 0.424 0.489 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.634 0.647 ;
        RECT MASK 1 -0.042 0.553 0.634 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.634 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.634 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.15 0.425 0.35 0.463 ;
      RECT MASK 1 0.316 0.155 0.35 0.425 ;
      RECT MASK 1 0.228 0.117 0.35 0.155 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.666 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.518 0.55 ;
      RECT 0.215 0.15 0.451 0.2 ;
      RECT 0.074 0.05 0.518 0.15 ;
    LAYER PO ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AO21B_0P5

MACRO SAEDRVT14_AOI21_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.444 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.222 0.202 0.414 ;
        RECT 0.168 0.222 0.202 0.414 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.199 0.128 0.377 ;
        RECT 0.094 0.199 0.128 0.377 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.199 0.276 0.377 ;
        RECT 0.242 0.199 0.276 0.377 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.316 0.146 0.35 0.415 ;
        RECT MASK 1 0.23 0.112 0.35 0.146 ;
        RECT 0.316 0.112 0.35 0.415 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.486 0.647 ;
        RECT MASK 1 -0.042 0.553 0.486 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.486 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.486 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.094 0.454 0.304 0.488 ;
      RECT MASK 1 0.094 0.417 0.128 0.454 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.518 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.37 0.55 ;
      RECT 0.229 0.35 0.37 0.4 ;
      RECT 0.155 0.2 0.289 0.25 ;
      RECT 0.074 0.15 0.289 0.2 ;
      RECT 0.074 0.05 0.37 0.15 ;
    LAYER PO ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AOI21_0P5

MACRO SAEDRVT14_OR2_MM_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.518 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.214 0.225 0.244 0.255 ;
      LAYER M2 ;
        RECT MASK 1 0.192 0.223 0.352 0.257 ;
        RECT 0.192 0.223 0.352 0.257 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.114 0.345 0.144 0.375 ;
      LAYER M2 ;
        RECT 0.011 0.343 0.17 0.377 ;
        RECT MASK 1 0.011 0.343 0.17 0.377 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.118 0.424 0.458 ;
        RECT 0.39 0.118 0.424 0.458 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.56 0.647 ;
        RECT MASK 1 -0.042 0.553 0.56 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.048 0.56 0.046 ;
        RECT MASK 1 -0.042 -0.048 0.56 0.046 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.226 0.454 0.35 0.488 ;
      RECT MASK 1 0.316 0.145 0.35 0.454 ;
      RECT MASK 1 0.15 0.111 0.35 0.145 ;
      RECT MASK 1 0.112 0.205 0.146 0.434 ;
      RECT MASK 1 0.212 0.205 0.246 0.389 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.592 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.444 0.55 ;
      RECT 0.155 0.4 0.303 0.45 ;
      RECT 0.074 0.05 0.444 0.15 ;
    LAYER PO ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OR2_MM_0P5

MACRO SAEDRVT14_NR3_0P75
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.74 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.199 0.276 0.418 ;
        RECT MASK 1 0.242 0.199 0.276 0.418 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.199 0.202 0.505 ;
        RECT MASK 1 0.168 0.199 0.202 0.505 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.212 0.128 0.441 ;
        RECT MASK 1 0.094 0.212 0.128 0.441 ;
    END
  END A3
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.101 0.646 0.472 ;
        RECT MASK 1 0.612 0.101 0.646 0.472 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.782 0.647 ;
        RECT MASK 1 -0.042 0.553 0.782 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.782 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.782 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.437 0.454 0.572 0.488 ;
      RECT MASK 1 0.538 0.146 0.572 0.454 ;
      RECT MASK 1 0.437 0.112 0.572 0.146 ;
      RECT MASK 1 0.316 0.316 0.35 0.488 ;
      RECT MASK 1 0.427 0.316 0.461 0.414 ;
      RECT MASK 1 0.316 0.282 0.461 0.316 ;
      RECT MASK 1 0.427 0.186 0.461 0.282 ;
      RECT MASK 1 0.316 0.146 0.35 0.282 ;
      RECT MASK 1 0.146 0.112 0.35 0.146 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.814 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.666 0.55 ;
      RECT 0.074 0.35 0.37 0.45 ;
      RECT 0.518 0.4 0.666 0.45 ;
      RECT 0.074 0.2 0.289 0.25 ;
      RECT 0.37 0.2 0.518 0.25 ;
      RECT 0.074 0.05 0.666 0.2 ;
    LAYER PO ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_NR3_0P75

MACRO SAEDRVT14_MUXI2_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.666 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.189 0.285 0.219 0.315 ;
      LAYER M2 ;
        RECT 0.182 0.283 0.438 0.317 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.464 0.176 0.498 0.424 ;
        RECT 0.464 0.176 0.498 0.424 ;
    END
  END D1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.353 0.225 0.383 0.255 ;
      LAYER M2 ;
        RECT 0.17 0.223 0.385 0.257 ;
        RECT MASK 1 0.17 0.223 0.385 0.257 ;
    END
  END S
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.538 0.102 0.572 0.498 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.046 0.553 0.708 0.647 ;
        RECT MASK 1 -0.046 0.553 0.708 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.046 -0.047 0.708 0.047 ;
        RECT MASK 1 -0.046 -0.047 0.708 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.351 0.176 0.385 0.424 ;
      RECT MASK 1 0.187 0.123 0.221 0.326 ;
    LAYER NWELL ;
      RECT -0.078 0.3 0.74 0.6 ;
    LAYER DIFF ;
      RECT 0.07 0.45 0.592 0.55 ;
      RECT 0.07 0.05 0.592 0.15 ;
    LAYER PO ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_MUXI2_U_0P5

MACRO SAEDRVT14_EO2_V1_0P75
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.74 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.244 0.285 0.274 0.315 ;
      LAYER M1 ;
        RECT MASK 1 0.242 0.215 0.276 0.365 ;
        RECT 0.242 0.215 0.276 0.365 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.102 0.128 0.484 ;
        RECT MASK 1 0.094 0.136 0.128 0.484 ;
        RECT MASK 1 0.612 0.136 0.646 0.339 ;
        RECT MASK 1 0.094 0.102 0.646 0.136 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.538 0.176 0.572 0.411 ;
        RECT MASK 1 0.464 0.377 0.572 0.411 ;
        RECT MASK 1 0.538 0.21 0.572 0.377 ;
        RECT MASK 1 0.371 0.176 0.572 0.21 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.782 0.647 ;
        RECT MASK 1 -0.042 0.553 0.782 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.782 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.782 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.39 0.464 0.646 0.498 ;
      RECT MASK 1 0.39 0.396 0.424 0.464 ;
      RECT MASK 1 0.612 0.379 0.646 0.464 ;
      RECT MASK 1 0.168 0.464 0.35 0.498 ;
      RECT MASK 1 0.168 0.176 0.202 0.464 ;
      RECT MASK 1 0.316 0.282 0.35 0.464 ;
      RECT MASK 1 0.39 0.267 0.498 0.317 ;
    LAYER VIA1 ;
      RECT 0.442 0.285 0.472 0.315 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.814 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.35 0.666 0.55 ;
      RECT 0.074 0.15 0.215 0.2 ;
      RECT 0.074 0.05 0.666 0.15 ;
    LAYER PO ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_EO2_V1_0P75

MACRO SAEDRVT14_NR4_0P75
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.814 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.339 0.345 0.369 0.375 ;
      LAYER M2 ;
        RECT 0.314 0.343 0.479 0.377 ;
        RECT MASK 1 0.314 0.343 0.479 0.377 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.265 0.465 0.295 0.495 ;
      LAYER M2 ;
        RECT 0.189 0.463 0.339 0.497 ;
        RECT MASK 1 0.189 0.463 0.339 0.497 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.2 0.202 0.464 ;
        RECT MASK 1 0.168 0.2 0.202 0.464 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.264 0.128 0.484 ;
        RECT MASK 1 0.094 0.264 0.128 0.484 ;
    END
  END A4
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.686 0.119 0.72 0.459 ;
        RECT 0.686 0.119 0.72 0.459 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.856 0.647 ;
        RECT MASK 1 -0.042 0.553 0.856 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.856 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.856 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.263 0.264 0.297 0.502 ;
      RECT MASK 1 0.52 0.443 0.623 0.488 ;
      RECT MASK 1 0.577 0.15 0.623 0.443 ;
      RECT MASK 1 0.52 0.112 0.623 0.15 ;
      RECT MASK 1 0.337 0.2 0.371 0.468 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.888 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.74 0.55 ;
      RECT 0.074 0.4 0.444 0.45 ;
      RECT 0.592 0.35 0.74 0.45 ;
      RECT 0.444 0.15 0.74 0.25 ;
      RECT 0.074 0.05 0.74 0.15 ;
    LAYER PO ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_NR4_0P75

MACRO SAEDRVT14_AN3_0P75
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.592 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.291 0.285 0.321 0.315 ;
      LAYER M2 ;
        RECT 0.237 0.283 0.385 0.317 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.213 0.345 0.243 0.375 ;
      LAYER M2 ;
        RECT 0.093 0.343 0.284 0.377 ;
        RECT MASK 1 0.093 0.343 0.284 0.377 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.112 0.128 0.378 ;
    END
  END A3
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.464 0.119 0.498 0.459 ;
        RECT MASK 1 0.464 0.119 0.498 0.459 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.634 0.647 ;
        RECT MASK 1 -0.042 0.553 0.634 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.634 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.634 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.15 0.45 0.432 0.488 ;
      RECT MASK 1 0.398 0.148 0.432 0.45 ;
      RECT MASK 1 0.304 0.114 0.432 0.148 ;
      RECT MASK 1 0.289 0.26 0.323 0.41 ;
      RECT MASK 1 0.211 0.259 0.245 0.409 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.666 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.511 0.55 ;
      RECT 0.377 0.35 0.511 0.4 ;
      RECT 0.289 0.2 0.377 0.25 ;
      RECT 0.074 0.05 0.511 0.2 ;
    LAYER PO ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AN3_0P75

MACRO SAEDRVT14_OAI311_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.962 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.234 0.35 0.418 ;
        RECT MASK 1 0.316 0.234 0.35 0.418 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.237 0.276 0.506 ;
        RECT MASK 1 0.242 0.237 0.276 0.506 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.24 0.128 0.458 ;
        RECT MASK 1 0.094 0.24 0.128 0.458 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.464 0.2 0.498 0.377 ;
        RECT 0.464 0.2 0.498 0.377 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.222 0.424 0.397 ;
        RECT 0.39 0.222 0.424 0.397 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.834 0.107 0.868 0.496 ;
        RECT MASK 1 0.834 0.107 0.868 0.496 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.004 0.647 ;
        RECT MASK 1 -0.042 0.553 1.004 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.004 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.004 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.684 0.319 0.722 0.496 ;
      RECT MASK 1 0.684 0.285 0.792 0.319 ;
      RECT MASK 1 0.684 0.107 0.722 0.285 ;
      RECT MASK 1 0.367 0.458 0.574 0.496 ;
      RECT MASK 1 0.536 0.319 0.574 0.458 ;
      RECT MASK 1 0.536 0.285 0.644 0.319 ;
      RECT MASK 1 0.536 0.107 0.574 0.285 ;
      RECT MASK 1 0.15 0.102 0.388 0.14 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.036 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.888 0.55 ;
      RECT 0.155 0.4 0.303 0.45 ;
      RECT 0.807 0.4 0.888 0.45 ;
      RECT 0.229 0.35 0.303 0.4 ;
      RECT 0.451 0.15 0.525 0.2 ;
      RECT 0.807 0.15 0.888 0.2 ;
      RECT 0.074 0.05 0.888 0.15 ;
    LAYER PO ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OAI311_1

MACRO SAEDRVT14_AN2_MM_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.518 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.186 0.202 0.412 ;
        RECT MASK 1 0.168 0.186 0.202 0.412 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.091 0.128 0.392 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 0.123 0.424 0.477 ;
        RECT MASK 1 0.39 0.123 0.424 0.477 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.56 0.647 ;
        RECT MASK 1 -0.042 0.553 0.56 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.56 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.56 0.047 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.3 0.592 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.444 0.55 ;
      RECT 0.074 0.15 0.296 0.2 ;
      RECT 0.074 0.05 0.444 0.15 ;
    LAYER PO ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AN2_MM_0P5

MACRO SAEDRVT14_AN2B_MM_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.666 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.192 0.424 0.408 ;
        RECT 0.39 0.192 0.424 0.408 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.163 0.128 0.435 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.536 0.144 0.574 0.498 ;
        RECT 0.536 0.144 0.574 0.498 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.049 0.553 0.708 0.647 ;
        RECT MASK 1 -0.049 0.553 0.708 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.708 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.708 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.168 0.324 0.202 0.477 ;
      RECT MASK 1 0.168 0.276 0.285 0.324 ;
      RECT MASK 1 0.168 0.123 0.202 0.276 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.74 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.592 0.55 ;
      RECT 0.222 0.35 0.592 0.4 ;
      RECT 0.222 0.2 0.592 0.25 ;
      RECT 0.074 0.05 0.592 0.2 ;
    LAYER PO ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AN2B_MM_1

MACRO SAEDRVT14_OA21_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.592 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.19 0.276 0.41 ;
        RECT MASK 1 0.242 0.19 0.276 0.41 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.115 0.465 0.145 0.495 ;
      LAYER M2 ;
        RECT -0.031 0.463 0.171 0.497 ;
        RECT MASK 1 -0.031 0.463 0.171 0.497 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.313 0.345 0.343 0.375 ;
      LAYER M2 ;
        RECT 0.243 0.343 0.43 0.377 ;
        RECT MASK 1 0.243 0.343 0.43 0.377 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.464 0.118 0.498 0.458 ;
        RECT MASK 1 0.464 0.118 0.498 0.458 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 0.553 0.634 0.647 ;
        RECT -0.042 0.553 0.634 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.634 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.634 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.107 0.288 0.153 0.506 ;
      RECT MASK 1 0.307 0.276 0.353 0.41 ;
      RECT MASK 1 0.093 0.112 0.31 0.15 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.666 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.518 0.55 ;
      RECT 0.37 0.35 0.518 0.4 ;
      RECT 0.37 0.2 0.518 0.25 ;
      RECT 0.074 0.15 0.155 0.2 ;
      RECT 0.289 0.15 0.518 0.2 ;
      RECT 0.074 0.05 0.518 0.15 ;
    LAYER PO ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OA21_1

MACRO SAEDRVT14_OR2_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.518 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.186 0.276 0.414 ;
        RECT 0.242 0.186 0.276 0.414 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.186 0.128 0.414 ;
        RECT 0.094 0.186 0.128 0.414 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.118 0.424 0.458 ;
        RECT 0.39 0.118 0.424 0.458 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.56 0.647 ;
        RECT MASK 1 -0.042 0.553 0.56 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.56 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.56 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.222 0.454 0.35 0.488 ;
      RECT MASK 1 0.316 0.146 0.35 0.454 ;
      RECT MASK 1 0.146 0.112 0.35 0.146 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.592 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.444 0.55 ;
      RECT 0.155 0.4 0.296 0.45 ;
      RECT 0.074 0.05 0.444 0.15 ;
    LAYER PO ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OR2_0P5

MACRO SAEDRVT14_AO33_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.888 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.393 0.225 0.423 0.255 ;
      LAYER M2 ;
        RECT MASK 1 0.234 0.223 0.431 0.257 ;
        RECT 0.234 0.223 0.431 0.257 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.505 0.285 0.535 0.315 ;
      LAYER M2 ;
        RECT 0.433 0.283 0.618 0.317 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.603 0.202 0.633 0.232 ;
      LAYER M2 ;
        RECT 0.599 0.2 0.796 0.234 ;
        RECT MASK 1 0.599 0.2 0.796 0.234 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.316 0.225 0.35 0.419 ;
        RECT 0.316 0.225 0.35 0.419 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.089 0.202 0.378 ;
        RECT MASK 1 0.168 0.089 0.202 0.378 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.159 0.128 0.419 ;
        RECT 0.094 0.159 0.128 0.419 ;
    END
  END B3
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.763 0.105 0.793 0.135 ;
      LAYER M2 ;
        RECT MASK 1 0.761 0.103 0.987 0.137 ;
        RECT 0.761 0.103 0.987 0.137 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.93 0.647 ;
        RECT MASK 1 -0.042 0.553 0.93 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.93 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.93 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.15 0.459 0.7 0.497 ;
      RECT MASK 1 0.761 0.089 0.795 0.489 ;
      RECT MASK 1 0.384 0.382 0.719 0.416 ;
      RECT MASK 1 0.685 0.155 0.719 0.382 ;
      RECT MASK 1 0.306 0.117 0.719 0.155 ;
      RECT MASK 1 0.599 0.2 0.645 0.342 ;
      RECT MASK 1 0.497 0.2 0.543 0.342 ;
      RECT MASK 1 0.385 0.2 0.431 0.342 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.962 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.814 0.55 ;
      RECT 0.303 0.15 0.585 0.2 ;
      RECT 0.074 0.05 0.814 0.15 ;
    LAYER PO ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AO33_U_0P5

MACRO SAEDRVT14_ND2_CDC_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.37 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.163 0.128 0.435 ;
        RECT MASK 1 0.094 0.163 0.128 0.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.274 0.276 0.477 ;
        RECT MASK 1 0.242 0.274 0.276 0.477 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.091 0.276 0.224 ;
        RECT MASK 1 0.168 0.224 0.202 0.509 ;
        RECT MASK 1 0.168 0.188 0.276 0.224 ;
        RECT MASK 1 0.242 0.091 0.276 0.188 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.55 0.412 0.647 ;
        RECT MASK 1 -0.042 0.55 0.412 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.412 0.05 ;
        RECT MASK 1 -0.042 -0.047 0.412 0.05 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.3 0.444 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.296 0.55 ;
      RECT 0.074 0.05 0.296 0.25 ;
    LAYER PO ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_ND2_CDC_1

MACRO SAEDRVT14_NR2_MM_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.37 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.16 0.276 0.363 ;
        RECT 0.242 0.16 0.276 0.363 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.159 0.128 0.383 ;
        RECT MASK 1 0.094 0.159 0.128 0.383 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.093 0.202 0.441 ;
        RECT MASK 1 0.236 0.441 0.27 0.509 ;
        RECT MASK 1 0.168 0.403 0.27 0.441 ;
        RECT MASK 1 0.168 0.093 0.202 0.403 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.412 0.647 ;
        RECT MASK 1 -0.042 0.553 0.412 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.412 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.412 0.047 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.299 0.444 0.619 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.296 0.55 ;
      RECT 0.074 0.05 0.296 0.15 ;
    LAYER PO ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_NR2_MM_0P5

MACRO SAEDRVT14_ND3_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.74 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.204 0.35 0.423 ;
        RECT MASK 1 0.316 0.204 0.35 0.423 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.103 0.276 0.419 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.111 0.128 0.444 ;
        RECT MASK 1 0.094 0.111 0.128 0.444 ;
    END
  END A3
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.119 0.646 0.497 ;
        RECT MASK 1 0.612 0.119 0.646 0.497 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.782 0.647 ;
        RECT MASK 1 -0.042 0.553 0.782 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.782 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.782 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.464 0.452 0.572 0.486 ;
      RECT MASK 1 0.538 0.149 0.572 0.452 ;
      RECT MASK 1 0.464 0.115 0.572 0.149 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.814 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.666 0.55 ;
      RECT 0.074 0.35 0.289 0.4 ;
      RECT 0.37 0.35 0.666 0.4 ;
      RECT 0.074 0.2 0.289 0.25 ;
      RECT 0.518 0.15 0.666 0.25 ;
      RECT 0.074 0.15 0.37 0.2 ;
      RECT 0.074 0.05 0.666 0.15 ;
    LAYER PO ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_ND3_0P5

MACRO SAEDRVT14_OAI31_0P75
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.814 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.177 0.276 0.356 ;
        RECT MASK 1 0.242 0.177 0.276 0.356 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.199 0.202 0.488 ;
        RECT 0.168 0.199 0.202 0.488 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.168 0.128 0.418 ;
        RECT 0.094 0.168 0.128 0.418 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.176 0.35 0.354 ;
        RECT MASK 1 0.316 0.176 0.35 0.354 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.686 0.119 0.72 0.459 ;
        RECT MASK 1 0.686 0.119 0.72 0.459 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.856 0.647 ;
        RECT MASK 1 -0.042 0.553 0.856 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.856 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.856 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.52 0.443 0.623 0.488 ;
      RECT MASK 1 0.577 0.15 0.623 0.443 ;
      RECT MASK 1 0.52 0.112 0.623 0.15 ;
      RECT MASK 1 0.312 0.422 0.424 0.46 ;
      RECT MASK 1 0.39 0.403 0.424 0.422 ;
      RECT MASK 1 0.39 0.369 0.517 0.403 ;
      RECT MASK 1 0.39 0.158 0.424 0.369 ;
      RECT MASK 1 0.483 0.192 0.517 0.369 ;
      RECT MASK 1 0.168 0.102 0.354 0.136 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.888 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.74 0.55 ;
      RECT 0.074 0.4 0.363 0.45 ;
      RECT 0.215 0.35 0.363 0.4 ;
      RECT 0.074 0.15 0.289 0.2 ;
      RECT 0.363 0.15 0.444 0.2 ;
      RECT 0.074 0.05 0.74 0.15 ;
    LAYER PO ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OAI31_0P75

MACRO SAEDRVT14_OAI222_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.184 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.538 0.226 0.572 0.437 ;
        RECT MASK 1 0.538 0.226 0.572 0.437 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.688 0.345 0.718 0.375 ;
      LAYER M2 ;
        RECT MASK 1 0.673 0.343 0.915 0.377 ;
        RECT 0.673 0.343 0.915 0.377 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.255 0.35 0.415 ;
        RECT MASK 1 0.316 0.255 0.35 0.415 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.429 0.285 0.459 0.315 ;
      LAYER M2 ;
        RECT 0.343 0.283 0.498 0.317 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.256 0.276 0.404 ;
        RECT MASK 1 0.242 0.256 0.276 0.404 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.199 0.128 0.488 ;
        RECT MASK 1 0.094 0.199 0.128 0.488 ;
    END
  END C2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 1.056 0.089 1.09 0.511 ;
        RECT 1.056 0.089 1.09 0.511 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.226 0.647 ;
        RECT MASK 1 -0.042 0.553 1.226 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.226 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.226 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.908 0.324 0.942 0.511 ;
      RECT MASK 1 0.908 0.283 1.016 0.324 ;
      RECT MASK 1 0.908 0.089 0.942 0.283 ;
      RECT MASK 1 0.213 0.464 0.81 0.498 ;
      RECT MASK 1 0.76 0.46 0.81 0.464 ;
      RECT MASK 1 0.76 0.324 0.796 0.46 ;
      RECT MASK 1 0.76 0.283 0.868 0.324 ;
      RECT MASK 1 0.76 0.14 0.794 0.283 ;
      RECT MASK 1 0.512 0.102 0.794 0.14 ;
      RECT MASK 1 0.683 0.259 0.723 0.412 ;
      RECT MASK 1 0.421 0.258 0.467 0.411 ;
      RECT MASK 1 0.304 0.166 0.7 0.2 ;
      RECT MASK 1 0.15 0.102 0.46 0.14 ;
      RECT 0.76 0.102 0.794 0.498 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.258 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 1.11 0.55 ;
      RECT 0.074 0.4 0.377 0.45 ;
      RECT 0.585 0.4 0.659 0.45 ;
      RECT 0.821 0.4 0.895 0.45 ;
      RECT 0.733 0.2 0.814 0.25 ;
      RECT 0.074 0.15 0.215 0.25 ;
      RECT 0.363 0.15 0.814 0.2 ;
      RECT 0.074 0.05 1.11 0.15 ;
    LAYER PO ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OAI222_0P5

MACRO SAEDRVT14_AOI311_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.962 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.158 0.35 0.418 ;
        RECT MASK 1 0.316 0.158 0.35 0.418 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.205 0.105 0.235 0.135 ;
      LAYER M2 ;
        RECT MASK 1 0.135 0.103 0.316 0.137 ;
        RECT 0.135 0.103 0.316 0.137 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.118 0.128 0.418 ;
        RECT MASK 1 0.094 0.118 0.128 0.418 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.464 0.199 0.498 0.436 ;
        RECT 0.464 0.199 0.498 0.436 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 0.199 0.424 0.405 ;
        RECT MASK 1 0.39 0.199 0.424 0.405 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.834 0.118 0.868 0.511 ;
        RECT 0.834 0.118 0.868 0.511 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.004 0.647 ;
        RECT MASK 1 -0.042 0.553 1.004 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.004 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.004 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.15 0.458 0.388 0.496 ;
      RECT MASK 1 0.684 0.321 0.722 0.488 ;
      RECT MASK 1 0.684 0.283 0.793 0.321 ;
      RECT MASK 1 0.684 0.118 0.722 0.283 ;
      RECT MASK 1 0.536 0.321 0.574 0.488 ;
      RECT MASK 1 0.536 0.283 0.644 0.321 ;
      RECT MASK 1 0.536 0.14 0.574 0.283 ;
      RECT MASK 1 0.38 0.102 0.574 0.14 ;
      RECT MASK 1 0.203 0.088 0.237 0.377 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.036 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.888 0.55 ;
      RECT 0.074 0.4 0.155 0.45 ;
      RECT 0.377 0.35 0.451 0.45 ;
      RECT 0.599 0.4 0.673 0.45 ;
      RECT 0.229 0.15 0.303 0.2 ;
      RECT 0.074 0.05 0.888 0.15 ;
    LAYER PO ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AOI311_0P5

MACRO SAEDRVT14_OA22_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.666 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.199 0.276 0.377 ;
        RECT 0.242 0.199 0.276 0.377 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.199 0.424 0.377 ;
        RECT 0.39 0.199 0.424 0.377 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.228 0.202 0.422 ;
        RECT MASK 1 0.168 0.228 0.202 0.422 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.263 0.128 0.488 ;
        RECT MASK 1 0.094 0.263 0.128 0.488 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.538 0.088 0.572 0.488 ;
        RECT MASK 1 0.538 0.088 0.572 0.488 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.708 0.647 ;
        RECT MASK 1 -0.042 0.553 0.708 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.708 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.708 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.242 0.444 0.498 0.482 ;
      RECT MASK 1 0.316 0.19 0.35 0.444 ;
      RECT MASK 1 0.464 0.246 0.498 0.444 ;
      RECT MASK 1 0.093 0.14 0.131 0.177 ;
      RECT MASK 1 0.093 0.102 0.431 0.14 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.74 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.592 0.55 ;
      RECT 0.155 0.4 0.229 0.45 ;
      RECT 0.074 0.05 0.592 0.15 ;
    LAYER PO ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OA22_U_0P5

MACRO SAEDRVT14_AN4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.666 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 0.19 0.424 0.41 ;
        RECT MASK 1 0.39 0.19 0.424 0.41 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.112 0.35 0.377 ;
        RECT MASK 1 0.316 0.112 0.35 0.377 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.165 0.276 0.41 ;
        RECT MASK 1 0.242 0.165 0.276 0.41 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.112 0.202 0.377 ;
        RECT MASK 1 0.168 0.112 0.202 0.377 ;
    END
  END A4
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.538 0.118 0.572 0.458 ;
        RECT 0.538 0.118 0.572 0.458 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.708 0.647 ;
        RECT MASK 1 -0.042 0.553 0.708 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.708 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.708 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.148 0.45 0.497 0.488 ;
      RECT MASK 1 0.463 0.15 0.497 0.45 ;
      RECT MASK 1 0.38 0.112 0.497 0.15 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.74 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.592 0.55 ;
      RECT 0.074 0.4 0.155 0.45 ;
      RECT 0.444 0.35 0.592 0.45 ;
      RECT 0.073 0.05 0.592 0.2 ;
    LAYER PO ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AN4_1

MACRO SAEDRVT14_NR3_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.74 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.212 0.276 0.45 ;
        RECT 0.242 0.212 0.276 0.45 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.199 0.202 0.511 ;
        RECT MASK 1 0.168 0.199 0.202 0.511 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.203 0.128 0.448 ;
        RECT MASK 1 0.094 0.203 0.128 0.448 ;
    END
  END A3
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.612 0.097 0.646 0.472 ;
        RECT 0.612 0.097 0.646 0.472 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.782 0.647 ;
        RECT MASK 1 -0.042 0.553 0.782 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.782 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.782 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.437 0.454 0.572 0.488 ;
      RECT MASK 1 0.538 0.146 0.572 0.454 ;
      RECT MASK 1 0.437 0.112 0.572 0.146 ;
      RECT MASK 1 0.316 0.316 0.35 0.488 ;
      RECT MASK 1 0.427 0.316 0.461 0.414 ;
      RECT MASK 1 0.316 0.282 0.461 0.316 ;
      RECT MASK 1 0.427 0.186 0.461 0.282 ;
      RECT MASK 1 0.316 0.146 0.35 0.282 ;
      RECT MASK 1 0.146 0.112 0.35 0.146 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.814 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.666 0.55 ;
      RECT 0.074 0.4 0.37 0.45 ;
      RECT 0.37 0.15 0.518 0.25 ;
      RECT 0.074 0.15 0.289 0.2 ;
      RECT 0.074 0.05 0.666 0.15 ;
    LAYER PO ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_NR3_0P5

MACRO SAEDRVT14_OAI21_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.444 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.221 0.202 0.413 ;
        RECT 0.168 0.221 0.202 0.413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.237 0.128 0.462 ;
        RECT 0.094 0.237 0.128 0.462 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.199 0.276 0.377 ;
        RECT 0.242 0.199 0.276 0.377 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.24 0.426 0.35 0.46 ;
        RECT MASK 1 0.316 0.187 0.35 0.426 ;
        RECT 0.316 0.187 0.35 0.46 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.486 0.647 ;
        RECT MASK 1 -0.042 0.553 0.486 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.486 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.486 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.094 0.136 0.128 0.182 ;
      RECT MASK 1 0.094 0.102 0.294 0.136 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.518 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.37 0.55 ;
      RECT 0.074 0.35 0.289 0.45 ;
      RECT 0.074 0.2 0.215 0.25 ;
      RECT 0.074 0.05 0.37 0.2 ;
    LAYER PO ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OAI21_0P5

MACRO SAEDRVT14_AOI22_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.814 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.199 0.276 0.377 ;
        RECT 0.242 0.199 0.276 0.377 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.088 0.424 0.313 ;
        RECT 0.39 0.088 0.424 0.313 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.222 0.202 0.418 ;
        RECT MASK 1 0.168 0.222 0.202 0.418 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.102 0.128 0.313 ;
        RECT 0.094 0.102 0.128 0.313 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.686 0.119 0.72 0.459 ;
        RECT MASK 1 0.686 0.119 0.72 0.459 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.856 0.647 ;
        RECT MASK 1 -0.042 0.553 0.856 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.856 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.856 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.094 0.458 0.426 0.496 ;
      RECT MASK 1 0.094 0.394 0.128 0.458 ;
      RECT MASK 1 0.52 0.443 0.623 0.488 ;
      RECT MASK 1 0.577 0.15 0.623 0.443 ;
      RECT MASK 1 0.52 0.112 0.623 0.15 ;
      RECT MASK 1 0.316 0.369 0.517 0.403 ;
      RECT MASK 1 0.483 0.192 0.517 0.369 ;
      RECT MASK 1 0.316 0.154 0.35 0.369 ;
      RECT MASK 1 0.226 0.116 0.35 0.154 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.888 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.74 0.55 ;
      RECT 0.363 0.4 0.444 0.45 ;
      RECT 0.155 0.15 0.289 0.2 ;
      RECT 0.074 0.05 0.74 0.15 ;
    LAYER PO ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AOI22_0P5

MACRO SAEDRVT14_INV_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.296 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.159 0.128 0.419 ;
        RECT 0.094 0.159 0.128 0.419 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.089 0.202 0.489 ;
        RECT 0.168 0.089 0.202 0.489 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 0.553 0.338 0.647 ;
        RECT -0.042 0.553 0.338 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 -0.048 0.338 0.046 ;
        RECT -0.042 -0.048 0.338 0.046 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.3 0.37 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.222 0.5 ;
      RECT 0.074 0.05 0.222 0.15 ;
    LAYER PO ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_INV_0P5

MACRO SAEDRVT14_OAI31_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.814 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.177 0.276 0.356 ;
        RECT 0.242 0.177 0.276 0.356 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.199 0.202 0.488 ;
        RECT MASK 1 0.168 0.199 0.202 0.488 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.168 0.128 0.418 ;
        RECT MASK 1 0.094 0.168 0.128 0.418 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.316 0.176 0.35 0.354 ;
        RECT 0.316 0.176 0.35 0.354 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.686 0.119 0.72 0.459 ;
        RECT MASK 1 0.686 0.119 0.72 0.459 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.856 0.647 ;
        RECT MASK 1 -0.042 0.553 0.856 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.856 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.856 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.52 0.443 0.623 0.488 ;
      RECT MASK 1 0.577 0.15 0.623 0.443 ;
      RECT MASK 1 0.52 0.112 0.623 0.15 ;
      RECT MASK 1 0.312 0.422 0.424 0.46 ;
      RECT MASK 1 0.39 0.403 0.424 0.422 ;
      RECT MASK 1 0.39 0.369 0.517 0.403 ;
      RECT MASK 1 0.39 0.158 0.424 0.369 ;
      RECT MASK 1 0.483 0.192 0.517 0.369 ;
      RECT MASK 1 0.168 0.102 0.354 0.136 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.888 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.74 0.55 ;
      RECT 0.074 0.4 0.363 0.45 ;
      RECT 0.289 0.35 0.363 0.4 ;
      RECT 0.074 0.15 0.215 0.2 ;
      RECT 0.363 0.15 0.444 0.2 ;
      RECT 0.074 0.05 0.74 0.15 ;
    LAYER PO ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OAI31_0P5

MACRO SAEDRVT14_OA33_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.888 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 0.262 0.424 0.414 ;
        RECT MASK 1 0.39 0.262 0.424 0.414 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.464 0.262 0.498 0.414 ;
        RECT 0.464 0.262 0.498 0.414 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.614 0.345 0.644 0.375 ;
      LAYER M2 ;
        RECT MASK 1 0.588 0.343 0.751 0.377 ;
        RECT 0.588 0.343 0.751 0.377 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.281 0.225 0.311 0.255 ;
      LAYER M2 ;
        RECT MASK 1 0.16 0.223 0.396 0.257 ;
        RECT 0.16 0.223 0.396 0.257 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.204 0.202 0.505 ;
        RECT MASK 1 0.168 0.204 0.202 0.505 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.186 0.128 0.458 ;
        RECT 0.094 0.186 0.128 0.458 ;
    END
  END B3
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.76 0.088 0.794 0.504 ;
        RECT 0.76 0.088 0.794 0.504 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.93 0.647 ;
        RECT MASK 1 -0.042 0.553 0.93 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.93 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.93 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.294 0.454 0.72 0.488 ;
      RECT MASK 1 0.686 0.222 0.72 0.454 ;
      RECT MASK 1 0.368 0.186 0.72 0.222 ;
      RECT MASK 1 0.606 0.262 0.652 0.414 ;
      RECT MASK 1 0.279 0.186 0.313 0.388 ;
      RECT MASK 1 0.146 0.112 0.668 0.146 ;
    LAYER NWELL ;
      RECT -0.074 0.299 0.962 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.814 0.55 ;
      RECT 0.155 0.4 0.437 0.45 ;
      RECT 0.525 0.15 0.673 0.2 ;
      RECT 0.074 0.05 0.814 0.15 ;
    LAYER PO ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OA33_U_0P5

MACRO SAEDRVT14_EO4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.072 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.289 0.345 0.319 0.375 ;
        RECT 0.54 0.345 0.57 0.375 ;
      LAYER M2 ;
        RECT MASK 1 0.264 0.343 0.602 0.377 ;
        RECT 0.264 0.343 0.602 0.377 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.176 0.128 0.333 ;
        RECT MASK 1 0.094 0.176 0.128 0.333 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.354 0.285 1.384 0.315 ;
        RECT 1.635 0.285 1.665 0.315 ;
      LAYER M2 ;
        RECT 1.336 0.283 1.691 0.317 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.798 0.225 1.828 0.255 ;
      LAYER M2 ;
        RECT 1.694 0.223 1.925 0.257 ;
        RECT MASK 1 1.694 0.223 1.925 0.257 ;
    END
  END A4
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 1.944 0.088 1.978 0.488 ;
        RECT 1.944 0.088 1.978 0.488 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 2.114 0.647 ;
        RECT MASK 1 -0.042 0.553 2.114 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 2.114 0.047 ;
        RECT MASK 1 -0.042 -0.047 2.114 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 1.204 0.464 1.73 0.498 ;
      RECT MASK 1 1.204 0.136 1.238 0.464 ;
      RECT MASK 1 1.204 0.102 1.632 0.136 ;
      RECT MASK 1 0.194 0.464 0.942 0.498 ;
      RECT MASK 1 0.686 0.136 0.72 0.464 ;
      RECT MASK 1 0.278 0.102 1.11 0.136 ;
      RECT MASK 1 1.056 0.283 1.09 0.488 ;
      RECT MASK 1 0.982 0.176 1.016 0.457 ;
      RECT MASK 1 1.87 0.176 1.904 0.45 ;
      RECT MASK 1 0.76 0.39 0.887 0.424 ;
      RECT MASK 1 0.76 0.197 0.794 0.39 ;
      RECT MASK 1 0.76 0.163 0.891 0.197 ;
      RECT MASK 1 1.633 0.176 1.667 0.418 ;
      RECT MASK 1 1.439 0.163 1.473 0.418 ;
      RECT MASK 1 1.278 0.176 1.312 0.418 ;
      RECT MASK 1 1.13 0.176 1.164 0.418 ;
      RECT MASK 1 0.612 0.176 0.646 0.418 ;
      RECT MASK 1 0.538 0.199 0.572 0.418 ;
      RECT MASK 1 0.287 0.199 0.321 0.418 ;
      RECT MASK 1 1.716 0.361 1.776 0.395 ;
      RECT MASK 1 1.716 0.136 1.75 0.361 ;
      RECT MASK 1 1.716 0.102 1.78 0.136 ;
      RECT MASK 1 0.146 0.361 0.237 0.395 ;
      RECT MASK 1 0.203 0.136 0.237 0.361 ;
      RECT MASK 1 0.146 0.102 0.237 0.136 ;
      RECT MASK 1 1.541 0.199 1.575 0.377 ;
      RECT MASK 1 1.352 0.199 1.386 0.377 ;
      RECT MASK 1 0.443 0.199 0.477 0.377 ;
      RECT MASK 1 0.365 0.199 0.399 0.377 ;
      RECT MASK 1 0.852 0.223 0.902 0.35 ;
      RECT MASK 1 1.796 0.176 1.83 0.325 ;
    LAYER M2 ;
      RECT MASK 1 0.968 0.343 1.924 0.377 ;
      RECT MASK 1 1.261 0.223 1.613 0.257 ;
      RECT MASK 1 0.835 0.223 1.172 0.257 ;
      RECT MASK 1 0.342 0.223 0.655 0.257 ;
    LAYER VIA1 ;
      RECT 1.872 0.345 1.902 0.375 ;
      RECT 0.984 0.345 1.014 0.375 ;
      RECT 1.058 0.285 1.088 0.315 ;
      RECT 0.762 0.285 0.792 0.315 ;
      RECT 0.445 0.285 0.475 0.315 ;
      RECT 0.205 0.285 0.235 0.315 ;
      RECT 1.543 0.225 1.573 0.255 ;
      RECT 1.28 0.225 1.31 0.255 ;
      RECT 1.132 0.225 1.162 0.255 ;
      RECT 0.86 0.225 0.89 0.255 ;
      RECT 0.614 0.225 0.644 0.255 ;
      RECT 0.367 0.225 0.397 0.255 ;
      RECT 1.718 0.165 1.748 0.195 ;
      RECT 1.441 0.165 1.471 0.195 ;
    LAYER NWELL ;
      RECT -0.074 0.3 2.146 0.6 ;
    LAYER DIFF ;
      RECT 0.888 0.45 1.998 0.55 ;
      RECT 1.554 0.4 1.998 0.45 ;
      RECT 1.85 0.35 1.998 0.4 ;
      RECT 0.074 0.45 0.814 0.55 ;
      RECT 0.074 0.4 0.37 0.45 ;
      RECT 0.518 0.4 0.814 0.45 ;
      RECT 1.85 0.2 1.998 0.25 ;
      RECT 0.888 0.15 1.11 0.2 ;
      RECT 1.702 0.15 1.998 0.2 ;
      RECT 0.888 0.05 1.998 0.15 ;
      RECT 0.074 0.15 0.222 0.2 ;
      RECT 0.666 0.15 0.814 0.2 ;
      RECT 0.074 0.05 0.814 0.15 ;
    LAYER PO ;
      RECT 2.065 0 2.079 0.6 ;
      RECT 1.991 0 2.005 0.6 ;
      RECT 1.917 0 1.931 0.6 ;
      RECT 1.843 0 1.857 0.6 ;
      RECT 1.769 0 1.783 0.6 ;
      RECT 1.695 0 1.709 0.6 ;
      RECT 1.621 0 1.635 0.6 ;
      RECT 1.547 0 1.561 0.6 ;
      RECT 1.473 0 1.487 0.6 ;
      RECT 1.399 0 1.413 0.6 ;
      RECT 1.325 0 1.339 0.6 ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_EO4_1

MACRO SAEDRVT14_MUX2_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.74 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.164 0.123 0.198 0.326 ;
        RECT MASK 1 0.164 0.123 0.198 0.326 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.46 0.176 0.494 0.424 ;
        RECT MASK 1 0.46 0.176 0.494 0.424 ;
    END
  END D1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.386 0.176 0.42 0.424 ;
        RECT MASK 1 0.386 0.176 0.42 0.424 ;
    END
  END S
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.608 0.123 0.642 0.477 ;
        RECT MASK 1 0.608 0.123 0.642 0.477 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.786 0.647 ;
        RECT MASK 1 -0.042 0.553 0.786 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.041 -0.047 0.786 0.047 ;
        RECT MASK 1 -0.041 -0.047 0.786 0.047 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.3 0.818 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.67 0.55 ;
      RECT 0.074 0.05 0.67 0.15 ;
    LAYER PO ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_MUX2_U_0P5

MACRO SAEDRVT14_OAI21_0P75
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.444 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.221 0.202 0.413 ;
        RECT 0.168 0.221 0.202 0.413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.237 0.128 0.462 ;
        RECT 0.094 0.237 0.128 0.462 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.199 0.276 0.377 ;
        RECT 0.242 0.199 0.276 0.377 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.24 0.426 0.35 0.46 ;
        RECT MASK 1 0.316 0.187 0.35 0.426 ;
        RECT 0.316 0.187 0.35 0.46 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.486 0.647 ;
        RECT MASK 1 -0.042 0.553 0.486 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.486 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.486 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.094 0.136 0.128 0.182 ;
      RECT MASK 1 0.094 0.102 0.294 0.136 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.518 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.37 0.55 ;
      RECT 0.074 0.35 0.289 0.45 ;
      RECT 0.074 0.2 0.215 0.25 ;
      RECT 0.074 0.05 0.37 0.2 ;
    LAYER PO ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OAI21_0P75

MACRO SAEDRVT14_AO222_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.258 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.834 0.19 0.868 0.344 ;
        RECT 0.834 0.19 0.868 0.344 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.984 0.285 1.014 0.315 ;
      LAYER M2 ;
        RECT 0.942 0.283 1.131 0.317 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.688 0.225 0.718 0.255 ;
      LAYER M2 ;
        RECT MASK 1 0.638 0.223 0.79 0.257 ;
        RECT 0.638 0.223 0.79 0.257 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.464 0.176 0.498 0.438 ;
        RECT 0.464 0.176 0.498 0.438 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.186 0.35 0.364 ;
        RECT MASK 1 0.316 0.186 0.35 0.364 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.106 0.128 0.482 ;
        RECT MASK 1 0.094 0.106 0.128 0.482 ;
    END
  END C2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.13 0.096 1.164 0.493 ;
        RECT MASK 1 1.13 0.096 1.164 0.493 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.3 0.647 ;
        RECT MASK 1 -0.042 0.553 1.3 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.3 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.3 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.39 0.464 0.646 0.498 ;
      RECT MASK 1 0.39 0.424 0.424 0.464 ;
      RECT MASK 1 0.168 0.39 0.424 0.424 ;
      RECT MASK 1 0.686 0.461 0.942 0.495 ;
      RECT MASK 1 0.686 0.421 0.72 0.461 ;
      RECT MASK 1 0.538 0.387 0.72 0.421 ;
      RECT MASK 1 0.76 0.384 1.09 0.418 ;
      RECT MASK 1 0.76 0.15 0.794 0.384 ;
      RECT MASK 1 1.056 0.117 1.09 0.384 ;
      RECT MASK 1 0.39 0.116 0.794 0.15 ;
      RECT MASK 1 0.982 0.19 1.016 0.344 ;
      RECT MASK 1 0.686 0.19 0.72 0.344 ;
      RECT MASK 1 0.538 0.21 0.646 0.258 ;
      RECT MASK 1 0.168 0.146 0.202 0.199 ;
      RECT MASK 1 0.168 0.112 0.35 0.146 ;
      RECT MASK 1 0.834 0.116 0.989 0.15 ;
      RECT 0.686 0.19 0.72 0.344 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.332 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 1.184 0.55 ;
      RECT 0.074 0.4 0.74 0.45 ;
      RECT 1.036 0.35 1.184 0.45 ;
      RECT 0.296 0.35 0.592 0.4 ;
      RECT 0.296 0.2 0.444 0.25 ;
      RECT 0.592 0.2 0.74 0.25 ;
      RECT 1.036 0.15 1.184 0.25 ;
      RECT 0.296 0.15 0.74 0.2 ;
      RECT 0.296 0.05 1.184 0.15 ;
      RECT 0.074 0.05 0.222 0.25 ;
    LAYER PO ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AO222_1

MACRO SAEDRVT14_EN3_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.406 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.772 0.405 0.802 0.435 ;
      LAYER M2 ;
        RECT 0.747 0.403 1.086 0.437 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.357 0.285 0.387 0.315 ;
      LAYER M2 ;
        RECT 0.345 0.283 0.679 0.317 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.265 0.128 0.42 ;
        RECT 0.094 0.265 0.128 0.42 ;
    END
  END A3
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 1.278 0.094 1.312 0.498 ;
        RECT 1.278 0.094 1.312 0.498 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.448 0.647 ;
        RECT MASK 1 -0.042 0.553 1.448 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.046 1.448 0.048 ;
        RECT MASK 1 -0.042 -0.046 1.448 0.048 ;
    END
  END VSS
  OBS
    LAYER M2 ;
      RECT MASK 1 0.814 0.343 1.158 0.377 ;
      RECT MASK 1 0.592 0.223 1.077 0.257 ;
      RECT MASK 1 0.18 0.223 0.511 0.257 ;
    LAYER VIA1 ;
      RECT 1.091 0.345 1.121 0.375 ;
      RECT 0.851 0.345 0.881 0.375 ;
      RECT 1.013 0.225 1.043 0.255 ;
      RECT 0.613 0.225 0.643 0.255 ;
      RECT 0.433 0.225 0.463 0.255 ;
      RECT 0.207 0.225 0.237 0.255 ;
      RECT 0.934 0.165 0.964 0.195 ;
      RECT 0.688 0.165 0.718 0.195 ;
      RECT 0.538 0.165 0.568 0.195 ;
      RECT 0.281 0.165 0.311 0.195 ;
    LAYER M1 ;
      RECT MASK 1 0.949 0.46 1.235 0.498 ;
      RECT MASK 1 1.201 0.137 1.235 0.46 ;
      RECT MASK 1 0.865 0.103 1.235 0.137 ;
      RECT MASK 1 0.849 0.211 0.883 0.498 ;
      RECT MASK 1 0.792 0.177 0.883 0.211 ;
      RECT MASK 1 0.15 0.46 0.239 0.498 ;
      RECT MASK 1 0.205 0.217 0.239 0.46 ;
      RECT MASK 1 0.15 0.183 0.239 0.217 ;
      RECT MASK 1 0.762 0.266 0.805 0.437 ;
      RECT MASK 1 0.932 0.163 0.967 0.42 ;
      RECT MASK 1 0.685 0.16 0.721 0.42 ;
      RECT MASK 1 0.534 0.163 0.571 0.42 ;
      RECT MASK 1 0.279 0.163 0.313 0.42 ;
      RECT MASK 1 1.089 0.177 1.123 0.379 ;
      RECT MASK 1 1.011 0.218 1.045 0.379 ;
      RECT MASK 1 0.431 0.178 0.465 0.379 ;
      RECT MASK 1 0.355 0.201 0.389 0.379 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.48 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 1.332 0.55 ;
      RECT 0.074 0.4 0.222 0.45 ;
      RECT 0.592 0.4 0.888 0.45 ;
      RECT 0.592 0.35 0.74 0.4 ;
      RECT 0.592 0.2 0.74 0.25 ;
      RECT 0.074 0.15 0.37 0.2 ;
      RECT 0.592 0.15 1.036 0.2 ;
      RECT 0.074 0.05 1.332 0.15 ;
    LAYER PO ;
      RECT 1.399 0 1.413 0.6 ;
      RECT 1.325 0 1.339 0.6 ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_EN3_U_0P5

MACRO SAEDRVT14_NR3B_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.888 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.162 0.128 0.448 ;
        RECT 0.094 0.162 0.128 0.448 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.199 0.35 0.384 ;
        RECT MASK 1 0.316 0.199 0.35 0.384 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.199 0.424 0.428 ;
        RECT 0.39 0.199 0.424 0.428 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.76 0.096 0.794 0.517 ;
        RECT 0.76 0.096 0.794 0.517 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.93 0.647 ;
        RECT MASK 1 -0.042 0.553 0.93 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.93 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.93 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.585 0.454 0.72 0.488 ;
      RECT MASK 1 0.686 0.146 0.72 0.454 ;
      RECT MASK 1 0.585 0.112 0.72 0.146 ;
      RECT MASK 1 0.226 0.454 0.498 0.488 ;
      RECT MASK 1 0.464 0.316 0.498 0.454 ;
      RECT MASK 1 0.575 0.316 0.609 0.414 ;
      RECT MASK 1 0.464 0.282 0.609 0.316 ;
      RECT MASK 1 0.575 0.186 0.609 0.282 ;
      RECT MASK 1 0.464 0.146 0.498 0.282 ;
      RECT MASK 1 0.315 0.112 0.498 0.146 ;
      RECT MASK 1 0.162 0.38 0.275 0.414 ;
      RECT MASK 1 0.241 0.184 0.275 0.38 ;
      RECT MASK 1 0.166 0.15 0.275 0.184 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.962 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.814 0.55 ;
      RECT 0.518 0.15 0.666 0.25 ;
      RECT 0.074 0.05 0.814 0.15 ;
    LAYER PO ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_NR3B_U_0P5

MACRO SAEDRVT14_AN2_MM_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.592 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.186 0.202 0.412 ;
        RECT MASK 1 0.168 0.186 0.202 0.412 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.127 0.128 0.392 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.464 0.15 0.498 0.441 ;
        RECT MASK 1 0.412 0.401 0.498 0.441 ;
        RECT MASK 1 0.464 0.19 0.498 0.401 ;
        RECT MASK 1 0.412 0.15 0.498 0.19 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.634 0.647 ;
        RECT MASK 1 -0.042 0.553 0.634 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.634 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.634 0.047 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.3 0.666 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.518 0.55 ;
      RECT 0.296 0.35 0.518 0.45 ;
      RECT 0.296 0.2 0.518 0.25 ;
      RECT 0.074 0.05 0.518 0.2 ;
    LAYER PO ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AN2_MM_2

MACRO SAEDRVT14_ADDH_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.11 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.254 0.225 0.284 0.255 ;
        RECT 0.654 0.225 0.684 0.255 ;
      LAYER M2 ;
        RECT 0.237 0.223 0.707 0.257 ;
        RECT MASK 1 0.237 0.223 0.707 0.257 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 0.163 0.424 0.431 ;
        RECT MASK 1 0.39 0.163 0.424 0.431 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.123 0.128 0.477 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.982 0.123 1.016 0.477 ;
        RECT 0.982 0.123 1.016 0.477 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 0.553 1.152 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.152 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.152 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.834 0.169 0.868 0.431 ;
      RECT MASK 1 0.56 0.169 0.594 0.431 ;
      RECT MASK 1 0.252 0.169 0.286 0.431 ;
      RECT MASK 1 0.723 0.194 0.757 0.423 ;
    LAYER M2 ;
      RECT MASK 1 0.555 0.343 0.89 0.377 ;
      RECT -0.042 0.553 1.152 0.647 ;
      RECT 0.094 0.123 0.128 0.477 ;
    LAYER VIA1 ;
      RECT 0.836 0.345 0.866 0.375 ;
      RECT 0.562 0.345 0.592 0.375 ;
      RECT 0.725 0.285 0.755 0.315 ;
      RECT 0.467 0.285 0.497 0.315 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.184 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 1.036 0.55 ;
      RECT 0.222 0.4 0.666 0.45 ;
      RECT 0.222 0.15 0.518 0.2 ;
      RECT 0.074 0.05 1.036 0.15 ;
    LAYER PO ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_ADDH_0P5

MACRO SAEDRVT14_BUF_1P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.518 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.186 0.202 0.414 ;
        RECT MASK 1 0.168 0.186 0.202 0.414 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.118 0.35 0.458 ;
        RECT MASK 1 0.316 0.118 0.35 0.458 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.56 0.647 ;
        RECT MASK 1 -0.042 0.553 0.56 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.56 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.56 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.146 0.454 0.276 0.488 ;
      RECT MASK 1 0.242 0.146 0.276 0.454 ;
      RECT MASK 1 0.146 0.112 0.276 0.146 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.592 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.444 0.55 ;
      RECT 0.074 0.05 0.444 0.2 ;
    LAYER PO ;
      RECT 0.512 0 0.526 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_BUF_1P5

MACRO SAEDRVT14_BUF_ECO_3
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.036 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.908 0.092 0.942 0.484 ;
        RECT MASK 1 0.908 0.092 0.942 0.484 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.614 0.225 0.644 0.255 ;
      LAYER M1 ;
        RECT 0.612 0.102 0.646 0.48 ;
        RECT MASK 1 0.612 0.43 0.71 0.48 ;
        RECT MASK 1 0.612 0.152 0.646 0.43 ;
        RECT MASK 1 0.612 0.102 0.71 0.152 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.043 0.553 1.078 0.647 ;
        RECT MASK 1 -0.043 0.553 1.078 0.647 ;
        RECT MASK 1 0.094 0.379 0.128 0.553 ;
        RECT MASK 1 0.316 0.379 0.35 0.553 ;
        RECT MASK 1 0.538 0.379 0.572 0.553 ;
        RECT MASK 1 0.834 0.409 0.868 0.553 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.078 0.047 ;
        RECT MASK 1 0.094 0.047 0.128 0.203 ;
        RECT MASK 1 0.316 0.047 0.35 0.203 ;
        RECT MASK 1 0.538 0.047 0.572 0.203 ;
        RECT MASK 1 0.834 0.047 0.868 0.165 ;
        RECT MASK 1 -0.042 -0.047 1.078 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.76 0.088 0.794 0.488 ;
      RECT MASK 1 0.4 0.43 0.498 0.48 ;
      RECT MASK 1 0.464 0.152 0.498 0.43 ;
      RECT MASK 1 0.4 0.102 0.498 0.152 ;
      RECT MASK 1 0.178 0.43 0.276 0.48 ;
      RECT MASK 1 0.242 0.152 0.276 0.43 ;
      RECT MASK 1 0.178 0.102 0.276 0.152 ;
      RECT MASK 1 0.686 0.202 0.72 0.374 ;
      RECT MASK 1 0.39 0.202 0.424 0.374 ;
      RECT MASK 1 0.168 0.202 0.202 0.374 ;
    LAYER VIA1 ;
      RECT 0.762 0.285 0.792 0.315 ;
      RECT 0.688 0.285 0.718 0.315 ;
      RECT 0.392 0.285 0.422 0.315 ;
      RECT 0.17 0.285 0.2 0.315 ;
      RECT 0.466 0.225 0.496 0.255 ;
      RECT 0.244 0.225 0.274 0.255 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.11 0.6 ;
    LAYER DIFF ;
      RECT 0.74 0.35 0.888 0.55 ;
      RECT 0.518 0.35 0.666 0.55 ;
      RECT 0.296 0.35 0.444 0.55 ;
      RECT 0.074 0.35 0.222 0.55 ;
      RECT 0.74 0.05 0.888 0.25 ;
      RECT 0.518 0.05 0.666 0.25 ;
      RECT 0.296 0.05 0.444 0.25 ;
      RECT 0.074 0.05 0.222 0.25 ;
    LAYER PO ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
    LAYER M2 ;
      RECT MASK 1 0.14 0.223 0.84 0.257 ;
  END
END SAEDRVT14_BUF_ECO_3

MACRO SAEDRVT14_BUF_S_1P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.518 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.201 0.128 0.388 ;
        RECT MASK 1 0.094 0.201 0.128 0.388 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.112 0.35 0.466 ;
        RECT MASK 1 0.297 0.41 0.35 0.466 ;
        RECT MASK 1 0.316 0.168 0.35 0.41 ;
        RECT MASK 1 0.297 0.112 0.35 0.168 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.56 0.647 ;
        RECT MASK 1 -0.042 0.553 0.56 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.56 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.56 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.205 0.256 0.283 0.322 ;
      RECT MASK 1 0.148 0.444 0.239 0.482 ;
      RECT MASK 1 0.205 0.322 0.239 0.444 ;
      RECT MASK 1 0.205 0.256 0.283 0.322 ;
      RECT MASK 1 0.205 0.151 0.239 0.256 ;
      RECT MASK 1 0.148 0.113 0.239 0.151 ;
    LAYER NWELL ;
      RECT -0.074 0.289 0.592 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.444 0.55 ;
      RECT 0.074 0.05 0.444 0.2 ;
    LAYER PO ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_BUF_S_1P5

MACRO SAEDRVT14_BUF_S_3
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.666 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.192 0.128 0.387 ;
        RECT MASK 1 0.094 0.192 0.128 0.387 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.402 0.405 0.432 0.435 ;
      LAYER M2 ;
        RECT 0.317 0.403 0.554 0.437 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.708 0.647 ;
        RECT MASK 1 -0.042 0.553 0.708 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.048 0.708 0.046 ;
        RECT MASK 1 -0.042 -0.048 0.708 0.046 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.148 0.448 0.239 0.486 ;
      RECT MASK 1 0.205 0.15 0.239 0.448 ;
      RECT MASK 1 0.148 0.112 0.239 0.15 ;
      RECT MASK 1 0.39 0.158 0.424 0.352 ;
    LAYER VIA1 ;
      RECT 0.392 0.165 0.422 0.195 ;
      RECT 0.207 0.165 0.237 0.195 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.74 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.35 0.592 0.55 ;
      RECT 0.074 0.05 0.592 0.25 ;
    LAYER PO ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_BUF_S_3

MACRO SAEDRVT14_BUF_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.444 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.211 0.202 0.364 ;
        RECT MASK 1 0.168 0.211 0.202 0.364 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.316 0.119 0.35 0.459 ;
        RECT 0.316 0.119 0.35 0.458 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.486 0.647 ;
        RECT MASK 1 -0.042 0.553 0.486 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.486 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.486 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.138 0.45 0.276 0.488 ;
      RECT MASK 1 0.242 0.146 0.276 0.45 ;
      RECT MASK 1 0.138 0.112 0.276 0.146 ;
    LAYER NWELL ;
      RECT -0.074 0.289 0.518 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.37 0.55 ;
      RECT 0.074 0.05 0.37 0.15 ;
    LAYER PO ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_BUF_U_0P5

MACRO SAEDRVT14_DEL_R2V1_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.518 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.163 0.202 0.435 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 0.102 0.424 0.498 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.56 0.647 ;
        RECT MASK 1 -0.042 0.553 0.56 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.56 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.56 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.233 0.464 0.35 0.498 ;
      RECT MASK 1 0.316 0.136 0.35 0.464 ;
      RECT MASK 1 0.232 0.102 0.35 0.136 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.592 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.444 0.55 ;
      RECT 0.296 0.35 0.444 0.45 ;
      RECT 0.296 0.15 0.444 0.25 ;
      RECT 0.074 0.05 0.444 0.15 ;
    LAYER PO ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_DEL_R2V1_1

MACRO SAEDRVT14_DEL_R2V2_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.814 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.131 0.158 0.165 0.418 ;
        RECT MASK 1 0.131 0.158 0.165 0.418 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.569 0.18 0.615 0.417 ;
        RECT MASK 1 0.512 0.383 0.615 0.417 ;
        RECT MASK 1 0.569 0.214 0.615 0.383 ;
        RECT MASK 1 0.512 0.18 0.615 0.214 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.856 0.647 ;
        RECT MASK 1 -0.042 0.553 0.856 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.856 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.856 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.316 0.458 0.72 0.496 ;
      RECT MASK 1 0.316 0.369 0.354 0.458 ;
      RECT MASK 1 0.685 0.369 0.72 0.458 ;
      RECT MASK 1 0.242 0.324 0.276 0.471 ;
      RECT MASK 1 0.242 0.278 0.439 0.324 ;
      RECT MASK 1 0.242 0.131 0.276 0.278 ;
      RECT MASK 1 0.316 0.14 0.354 0.229 ;
      RECT MASK 1 0.684 0.14 0.72 0.229 ;
      RECT MASK 1 0.316 0.102 0.72 0.14 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.888 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.35 0.74 0.55 ;
      RECT 0.074 0.05 0.74 0.25 ;
    LAYER PO ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_DEL_R2V2_2

MACRO SAEDRVT14_INV_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.518 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.244 0.165 0.274 0.195 ;
      LAYER M2 ;
        RECT 0.162 0.163 0.357 0.197 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.244 0.405 0.274 0.435 ;
      LAYER M2 ;
        RECT 0.162 0.403 0.356 0.437 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.56 0.647 ;
        RECT MASK 1 -0.042 0.553 0.56 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.56 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.56 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.149 0.403 0.351 0.469 ;
      RECT MASK 1 0.149 0.403 0.351 0.469 ;
      RECT MASK 1 0.159 0.082 0.202 0.403 ;
      RECT MASK 1 0.316 0.082 0.351 0.403 ;
      RECT MASK 1 0.242 0.158 0.276 0.329 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.592 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.35 0.444 0.55 ;
      RECT 0.074 0.05 0.444 0.25 ;
    LAYER PO ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_INV_4

MACRO SAEDRVT14_INV_S_1P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.37 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.159 0.128 0.419 ;
        RECT MASK 1 0.094 0.159 0.128 0.419 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.089 0.202 0.489 ;
        RECT MASK 1 0.168 0.089 0.202 0.489 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 0.553 0.412 0.647 ;
        RECT -0.042 0.553 0.412 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.412 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.412 0.047 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.3 0.444 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.296 0.55 ;
      RECT 0.074 0.05 0.296 0.2 ;
    LAYER PO ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_INV_S_1P5

MACRO SAEDRVT14_INV_S_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.37 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.159 0.128 0.419 ;
        RECT 0.094 0.159 0.128 0.419 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.089 0.202 0.489 ;
        RECT 0.168 0.089 0.202 0.489 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.412 0.647 ;
        RECT MASK 1 -0.042 0.553 0.412 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 -0.047 0.412 0.047 ;
        RECT -0.042 -0.047 0.412 0.047 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.3 0.444 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.35 0.296 0.55 ;
      RECT 0.074 0.05 0.296 0.25 ;
    LAYER PO ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_INV_S_2

MACRO SAEDRVT14_AOINV_IW_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.666 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.139 0.128 0.349 ;
        RECT MASK 1 0.094 0.139 0.128 0.349 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.368 0.276 0.402 ;
        RECT MASK 1 0.242 0.179 0.276 0.368 ;
        RECT MASK 1 0.168 0.145 0.276 0.179 ;
        RECT 0.242 0.145 0.276 0.402 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.708 0.647 ;
        RECT MASK 1 -0.042 0.553 0.708 0.647 ;
    END
  END VDD
  PIN VDDR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.102 0.466 0.132 0.496 ;
      LAYER M2 ;
        RECT -0.046 0.457 0.708 0.543 ;
        RECT MASK 1 -0.046 0.457 0.708 0.543 ;
    END
  END VDDR
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.708 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.708 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.094 0.464 0.196 0.498 ;
      RECT MASK 1 0.094 0.389 0.128 0.464 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.74 0.6 ;
    LAYER DIFF ;
      RECT 0.296 0.5 0.518 0.55 ;
      RECT 0.074 0.45 0.222 0.55 ;
      RECT 0.074 0.05 0.222 0.15 ;
      RECT 0.296 0.05 0.518 0.1 ;
    LAYER PO ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AOINV_IW_0P5

MACRO SAEDRVT14_AOINV_IW_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.666 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.139 0.128 0.349 ;
        RECT MASK 1 0.094 0.139 0.128 0.349 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.145 0.276 0.402 ;
        RECT MASK 1 0.168 0.368 0.276 0.402 ;
        RECT MASK 1 0.242 0.179 0.276 0.368 ;
        RECT MASK 1 0.168 0.145 0.276 0.179 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.708 0.647 ;
        RECT MASK 1 -0.042 0.553 0.708 0.647 ;
    END
  END VDD
  PIN VDDR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.102 0.466 0.132 0.496 ;
      LAYER M2 ;
        RECT -0.042 0.457 0.708 0.543 ;
        RECT MASK 1 -0.042 0.457 0.708 0.543 ;
    END
  END VDDR
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.708 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.708 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.094 0.464 0.196 0.498 ;
      RECT MASK 1 0.094 0.389 0.128 0.464 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.74 0.6 ;
    LAYER DIFF ;
      RECT 0.296 0.5 0.518 0.55 ;
      RECT 0.074 0.35 0.222 0.55 ;
      RECT 0.074 0.05 0.222 0.2 ;
      RECT 0.296 0.05 0.518 0.1 ;
    LAYER PO ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AOINV_IW_1

MACRO SAEDRVT14_AOINV_IW_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.74 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.139 0.128 0.349 ;
        RECT MASK 1 0.094 0.139 0.128 0.349 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.368 0.35 0.402 ;
        RECT MASK 1 0.316 0.179 0.35 0.368 ;
        RECT MASK 1 0.168 0.145 0.35 0.179 ;
        RECT 0.316 0.145 0.35 0.402 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.782 0.647 ;
        RECT MASK 1 -0.042 0.553 0.782 0.647 ;
    END
  END VDD
  PIN VDDR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.102 0.466 0.132 0.496 ;
        RECT 0.244 0.466 0.274 0.496 ;
      LAYER M2 ;
        RECT -0.042 0.457 0.782 0.543 ;
        RECT MASK 1 -0.042 0.457 0.782 0.543 ;
    END
  END VDDR
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.782 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.782 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.094 0.464 0.276 0.498 ;
      RECT MASK 1 0.094 0.389 0.128 0.464 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.814 0.6 ;
    LAYER DIFF ;
      RECT 0.37 0.5 0.592 0.55 ;
      RECT 0.074 0.35 0.296 0.55 ;
      RECT 0.074 0.05 0.296 0.2 ;
      RECT 0.37 0.05 0.592 0.1 ;
    LAYER PO ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AOINV_IW_2

MACRO SAEDRVT14_AOINV_IW_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.888 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.139 0.128 0.349 ;
        RECT MASK 1 0.094 0.139 0.128 0.349 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.464 0.145 0.498 0.402 ;
        RECT MASK 1 0.168 0.368 0.498 0.402 ;
        RECT MASK 1 0.464 0.179 0.498 0.368 ;
        RECT MASK 1 0.168 0.145 0.498 0.179 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.93 0.647 ;
        RECT MASK 1 -0.042 0.553 0.93 0.647 ;
    END
  END VDD
  PIN VDDR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.102 0.466 0.132 0.496 ;
        RECT 0.244 0.466 0.274 0.496 ;
        RECT 0.392 0.466 0.422 0.496 ;
      LAYER M2 ;
        RECT -0.042 0.457 0.93 0.543 ;
        RECT MASK 1 -0.042 0.457 0.93 0.543 ;
    END
  END VDDR
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.93 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.93 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.094 0.464 0.424 0.498 ;
      RECT MASK 1 0.094 0.389 0.128 0.464 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.962 0.6 ;
    LAYER DIFF ;
      RECT 0.518 0.5 0.74 0.55 ;
      RECT 0.074 0.35 0.444 0.55 ;
      RECT 0.074 0.05 0.444 0.2 ;
      RECT 0.518 0.05 0.74 0.1 ;
    LAYER PO ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AOINV_IW_4

MACRO SAEDRVT14_AOINV_IW_6
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.036 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.21 0.283 0.493 0.317 ;
        RECT MASK 1 0.21 0.283 0.493 0.317 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.368 0.646 0.402 ;
        RECT MASK 1 0.612 0.179 0.646 0.368 ;
        RECT MASK 1 0.168 0.145 0.646 0.179 ;
        RECT 0.612 0.145 0.646 0.402 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.079 0.647 ;
        RECT MASK 1 -0.042 0.553 1.078 0.647 ;
    END
  END VDD
  PIN VDDR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER VIA1 ;
        RECT 0.102 0.466 0.132 0.496 ;
        RECT 0.244 0.466 0.274 0.496 ;
        RECT 0.392 0.466 0.422 0.496 ;
        RECT 0.54 0.466 0.57 0.496 ;
      LAYER M2 ;
        RECT -0.042 0.457 1.078 0.543 ;
        RECT MASK 1 -0.042 0.457 1.078 0.543 ;
    END
  END VDDR
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.046 1.078 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.078 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.094 0.464 0.572 0.498 ;
      RECT MASK 1 0.094 0.389 0.128 0.464 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.11 0.6 ;
    LAYER DIFF ;
      RECT 0.666 0.5 0.888 0.55 ;
      RECT 0.074 0.35 0.592 0.55 ;
      RECT 0.074 0.05 0.592 0.2 ;
      RECT 0.666 0.05 0.888 0.1 ;
    LAYER PO ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AOINV_IW_6

MACRO SAEDRVT14_AN2_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.48 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.538 0.257 0.572 0.407 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.257 0.276 0.407 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.835 0.405 0.865 0.435 ;
        RECT 0.985 0.405 1.015 0.435 ;
        RECT 1.131 0.405 1.161 0.435 ;
      LAYER M2 ;
        RECT 0.824 0.403 1.324 0.437 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.554 1.526 0.648 ;
        RECT MASK 1 -0.042 0.554 1.526 0.648 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.526 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.526 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.146 0.439 0.763 0.479 ;
      RECT MASK 1 0.721 0.217 0.763 0.439 ;
      RECT MASK 1 0.442 0.181 0.763 0.217 ;
      RECT MASK 1 1.205 0.163 1.239 0.342 ;
      RECT MASK 1 1.057 0.163 1.091 0.342 ;
      RECT MASK 1 0.909 0.163 0.943 0.342 ;
    LAYER VIA1 ;
      RECT 1.207 0.185 1.237 0.215 ;
      RECT 1.059 0.185 1.089 0.215 ;
      RECT 0.911 0.185 0.941 0.215 ;
      RECT 0.724 0.185 0.754 0.215 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.558 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.35 1.41 0.55 ;
      RECT 0.074 0.2 0.74 0.25 ;
      RECT 0.074 0.05 1.41 0.2 ;
    LAYER PO ;
      RECT 1.473 0 1.487 0.6 ;
      RECT 1.399 0 1.413 0.6 ;
      RECT 1.325 0 1.339 0.6 ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AN2_8

MACRO SAEDRVT14_ND2_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.518 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.255 0.276 0.403 ;
        RECT 0.242 0.255 0.276 0.403 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.1 0.165 0.13 0.195 ;
      LAYER M2 ;
        RECT -0.001 0.163 0.183 0.197 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.304 0.225 0.334 0.255 ;
      LAYER M2 ;
        RECT 0.198 0.223 0.382 0.257 ;
        RECT MASK 1 0.198 0.223 0.382 0.257 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.56 0.647 ;
        RECT MASK 1 -0.042 0.553 0.56 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.56 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.56 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.161 0.444 0.399 0.478 ;
      RECT MASK 1 0.302 0.215 0.336 0.444 ;
      RECT MASK 1 0.238 0.181 0.336 0.215 ;
      RECT MASK 1 0.386 0.14 0.42 0.34 ;
      RECT MASK 1 0.098 0.14 0.132 0.336 ;
      RECT MASK 1 0.098 0.102 0.42 0.14 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.592 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.444 0.55 ;
      RECT 0.074 0.4 0.215 0.45 ;
      RECT 0.229 0.2 0.303 0.25 ;
      RECT 0.155 0.15 0.444 0.2 ;
      RECT 0.074 0.05 0.444 0.15 ;
    LAYER PO ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_ND2_0P5

MACRO SAEDRVT14_ND2_MM_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.518 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.316 0.261 0.35 0.477 ;
        RECT 0.316 0.261 0.35 0.477 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.166 0.202 0.456 ;
        RECT 0.168 0.166 0.202 0.456 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.178 0.276 0.509 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.56 0.647 ;
        RECT MASK 1 -0.042 0.553 0.56 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.56 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.56 0.047 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.3 0.593 0.6 ;
    LAYER DIFF ;
      RECT 0.148 0.35 0.371 0.55 ;
      RECT 0.074 0.05 0.444 0.25 ;
    LAYER PO ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_ND2_MM_1

MACRO SAEDRVT14_OA2BB2_V1_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.814 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.523 0.285 0.553 0.315 ;
      LAYER M2 ;
        RECT 0.437 0.283 0.747 0.317 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.627 0.225 0.657 0.255 ;
      LAYER M2 ;
        RECT 0.511 0.223 0.821 0.257 ;
        RECT MASK 1 0.511 0.223 0.821 0.257 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.205 0.202 0.488 ;
        RECT MASK 1 0.168 0.205 0.202 0.488 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.224 0.128 0.418 ;
        RECT MASK 1 0.094 0.224 0.128 0.418 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.449 0.345 0.479 0.375 ;
      LAYER M2 ;
        RECT 0.289 0.343 0.599 0.377 ;
        RECT MASK 1 0.289 0.343 0.599 0.377 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.861 0.647 ;
        RECT MASK 1 -0.042 0.553 0.861 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.861 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.861 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.462 0.458 0.669 0.496 ;
      RECT MASK 1 0.631 0.378 0.669 0.458 ;
      RECT MASK 1 0.331 0.395 0.369 0.488 ;
      RECT MASK 1 0.331 0.361 0.481 0.395 ;
      RECT MASK 1 0.447 0.14 0.481 0.361 ;
      RECT MASK 1 0.447 0.102 0.494 0.14 ;
      RECT MASK 1 0.257 0.214 0.397 0.28 ;
      RECT MASK 1 0.257 0.28 0.291 0.418 ;
      RECT MASK 1 0.257 0.214 0.397 0.28 ;
      RECT MASK 1 0.257 0.154 0.291 0.214 ;
      RECT MASK 1 0.15 0.116 0.291 0.154 ;
      RECT MASK 1 0.521 0.18 0.555 0.403 ;
      RECT MASK 1 0.619 0.18 0.665 0.329 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.893 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.74 0.55 ;
      RECT 0.074 0.05 0.666 0.15 ;
    LAYER PO ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OA2BB2_V1_0P5

MACRO SAEDRVT14_OA31_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.036 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.542 0.345 0.572 0.375 ;
      LAYER M2 ;
        RECT MASK 1 0.469 0.343 0.619 0.377 ;
        RECT 0.469 0.343 0.619 0.377 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.316 0.186 0.35 0.34 ;
        RECT 0.316 0.186 0.35 0.34 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.17 0.128 0.43 ;
        RECT 0.094 0.17 0.128 0.43 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.688 0.285 0.718 0.315 ;
      LAYER M2 ;
        RECT 0.646 0.283 0.796 0.317 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.908 0.117 0.942 0.493 ;
        RECT MASK 1 0.908 0.117 0.942 0.493 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.078 0.647 ;
        RECT MASK 1 -0.042 0.553 1.078 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.078 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.078 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.612 0.454 0.868 0.488 ;
      RECT MASK 1 0.834 0.143 0.868 0.454 ;
      RECT MASK 1 0.76 0.109 0.868 0.143 ;
      RECT MASK 1 0.39 0.454 0.572 0.488 ;
      RECT MASK 1 0.168 0.454 0.35 0.488 ;
      RECT MASK 1 0.316 0.414 0.35 0.454 ;
      RECT MASK 1 0.316 0.38 0.498 0.414 ;
      RECT MASK 1 0.686 0.237 0.72 0.414 ;
      RECT MASK 1 0.54 0.24 0.574 0.4 ;
      RECT MASK 1 0.168 0.112 0.72 0.146 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.11 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.962 0.55 ;
      RECT 0.074 0.4 0.666 0.45 ;
      RECT 0.814 0.4 0.962 0.45 ;
      RECT 0.518 0.35 0.666 0.4 ;
      RECT 0.666 0.2 0.814 0.25 ;
      RECT 0.666 0.15 0.962 0.2 ;
      RECT 0.518 0.05 0.962 0.15 ;
      RECT 0.074 0.05 0.222 0.25 ;
      RECT 0.296 0.05 0.444 0.2 ;
    LAYER PO ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OA31_U_0P5

MACRO SAEDRVT14_EN2_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.962 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.427 0.345 0.457 0.375 ;
      LAYER M2 ;
        RECT 0.407 0.343 0.647 0.377 ;
        RECT MASK 1 0.407 0.343 0.647 0.377 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.187 0.345 0.217 0.375 ;
      LAYER M2 ;
        RECT MASK 1 0.006 0.343 0.246 0.377 ;
        RECT 0.006 0.343 0.246 0.377 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.76 0.103 0.794 0.477 ;
        RECT 0.76 0.103 0.794 0.477 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.004 0.647 ;
        RECT MASK 1 -0.042 0.553 1.004 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.004 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.004 0.047 ;
    END
  END VSS
  OBS
    LAYER M2 ;
      RECT MASK 1 0.253 0.223 0.56 0.257 ;
    LAYER VIA1 ;
      RECT 0.505 0.225 0.535 0.255 ;
      RECT 0.277 0.225 0.307 0.255 ;
      RECT 0.615 0.165 0.645 0.195 ;
      RECT 0.353 0.165 0.383 0.195 ;
    LAYER M1 ;
      RECT MASK 1 0.608 0.163 0.65 0.416 ;
      RECT MASK 1 0.351 0.163 0.385 0.416 ;
      RECT MASK 1 0.181 0.274 0.223 0.416 ;
      RECT MASK 1 0.503 0.182 0.537 0.392 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.036 0.6 ;
    LAYER DIFF ;
      RECT 0.148 0.45 0.888 0.55 ;
      RECT 0.148 0.4 0.296 0.45 ;
      RECT 0.303 0.15 0.444 0.2 ;
      RECT 0.666 0.15 0.807 0.2 ;
      RECT 0.074 0.05 0.814 0.15 ;
    LAYER PO ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_EN2_0P5

MACRO SAEDRVT14_AOI222_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.184 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.577 0.225 0.607 0.255 ;
      LAYER M2 ;
        RECT 0.491 0.223 0.641 0.257 ;
        RECT MASK 1 0.491 0.223 0.641 0.257 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.688 0.285 0.718 0.315 ;
      LAYER M2 ;
        RECT 0.673 0.283 0.841 0.317 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.176 0.35 0.361 ;
        RECT MASK 1 0.316 0.176 0.35 0.361 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.464 0.173 0.498 0.36 ;
        RECT 0.464 0.173 0.498 0.36 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.199 0.276 0.387 ;
        RECT 0.242 0.199 0.276 0.387 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.11 0.128 0.377 ;
        RECT 0.094 0.11 0.128 0.377 ;
    END
  END C2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.056 0.118 1.09 0.458 ;
        RECT MASK 1 1.056 0.118 1.09 0.458 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.226 0.647 ;
        RECT MASK 1 -0.042 0.553 1.226 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.226 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.226 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.538 0.464 0.794 0.498 ;
      RECT MASK 1 0.76 0.365 0.794 0.464 ;
      RECT MASK 1 0.76 0.331 0.887 0.365 ;
      RECT MASK 1 0.853 0.191 0.887 0.331 ;
      RECT MASK 1 0.76 0.136 0.794 0.331 ;
      RECT MASK 1 0.228 0.102 0.794 0.136 ;
      RECT MASK 1 0.15 0.464 0.46 0.498 ;
      RECT MASK 1 0.89 0.442 0.993 0.487 ;
      RECT MASK 1 0.947 0.149 0.993 0.442 ;
      RECT MASK 1 0.89 0.111 0.993 0.149 ;
      RECT MASK 1 0.304 0.39 0.72 0.424 ;
      RECT MASK 1 0.681 0.199 0.725 0.35 ;
      RECT MASK 1 0.567 0.176 0.617 0.321 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.258 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 1.11 0.55 ;
      RECT 0.437 0.4 0.814 0.45 ;
      RECT 0.666 0.35 0.814 0.4 ;
      RECT 0.155 0.15 0.296 0.2 ;
      RECT 0.074 0.05 1.11 0.15 ;
    LAYER PO ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AOI222_0P5

MACRO SAEDRVT14_ND2_ECO_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.592 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.201 0.276 0.397 ;
        RECT MASK 1 0.242 0.201 0.276 0.397 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 0.201 0.424 0.397 ;
        RECT MASK 1 0.39 0.201 0.424 0.397 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.236 0.202 0.491 ;
        RECT MASK 1 0.168 0.439 0.378 0.491 ;
        RECT MASK 1 0.168 0.283 0.202 0.439 ;
        RECT MASK 1 0.094 0.236 0.202 0.283 ;
        RECT MASK 1 0.094 0.091 0.128 0.236 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.634 0.647 ;
        RECT MASK 1 -0.042 0.553 0.634 0.647 ;
        RECT MASK 1 0.094 0.364 0.128 0.553 ;
        RECT MASK 1 0.464 0.394 0.498 0.553 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.634 0.047 ;
        RECT MASK 1 0.464 0.047 0.498 0.206 ;
        RECT MASK 1 -0.042 -0.047 0.634 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.194 0.109 0.381 0.161 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.666 0.6 ;
    LAYER DIFF ;
      RECT 0.296 0.4 0.444 0.55 ;
      RECT 0.074 0.45 0.222 0.55 ;
      RECT 0.296 0.05 0.444 0.25 ;
      RECT 0.074 0.05 0.222 0.25 ;
    LAYER PO ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_ND2_ECO_1

MACRO SAEDRVT14_OA21_MM_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.666 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.213 0.405 0.243 0.435 ;
      LAYER M2 ;
        RECT 0.203 0.403 0.39 0.437 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.116 0.345 0.146 0.375 ;
      LAYER M2 ;
        RECT 0.021 0.343 0.19 0.377 ;
        RECT MASK 1 0.021 0.343 0.19 0.377 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 0.19 0.424 0.352 ;
        RECT MASK 1 0.39 0.19 0.424 0.352 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.538 0.112 0.572 0.501 ;
        RECT MASK 1 0.538 0.112 0.572 0.501 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.708 0.647 ;
        RECT MASK 1 -0.042 0.553 0.708 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.708 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.708 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.211 0.264 0.245 0.502 ;
      RECT MASK 1 0.107 0.247 0.153 0.418 ;
      RECT MASK 1 0.103 0.15 0.141 0.207 ;
      RECT MASK 1 0.103 0.112 0.388 0.15 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.74 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.592 0.55 ;
      RECT 0.444 0.35 0.592 0.4 ;
      RECT 0.074 0.2 0.222 0.25 ;
      RECT 0.444 0.2 0.592 0.25 ;
      RECT 0.074 0.05 0.592 0.2 ;
    LAYER PO ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OA21_MM_1

MACRO SAEDRVT14_OAI33_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.11 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.464 0.255 0.498 0.413 ;
        RECT MASK 1 0.464 0.255 0.498 0.413 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.538 0.255 0.572 0.413 ;
        RECT 0.538 0.255 0.572 0.413 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.658 0.345 0.688 0.375 ;
      LAYER M2 ;
        RECT 0.644 0.343 0.887 0.377 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.184 0.276 0.378 ;
        RECT MASK 1 0.242 0.184 0.276 0.378 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.199 0.202 0.447 ;
        RECT MASK 1 0.168 0.199 0.202 0.447 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.202 0.128 0.507 ;
        RECT 0.094 0.202 0.128 0.507 ;
    END
  END B3
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.982 0.089 1.016 0.511 ;
        RECT 0.982 0.089 1.016 0.511 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.152 0.647 ;
        RECT MASK 1 -0.042 0.553 1.152 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.152 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.152 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.834 0.319 0.868 0.511 ;
      RECT MASK 1 0.834 0.283 0.942 0.319 ;
      RECT MASK 1 0.834 0.089 0.868 0.283 ;
      RECT MASK 1 0.536 0.439 0.657 0.498 ;
      RECT MASK 1 0.308 0.439 0.429 0.473 ;
      RECT MASK 1 0.351 0.215 0.387 0.439 ;
      RECT MASK 1 0.76 0.215 0.794 0.419 ;
      RECT MASK 1 0.351 0.181 0.794 0.215 ;
      RECT MASK 1 0.653 0.257 0.693 0.397 ;
      RECT MASK 1 0.166 0.103 0.722 0.141 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.184 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 1.036 0.55 ;
      RECT 0.074 0.4 0.363 0.45 ;
      RECT 0.451 0.4 0.74 0.45 ;
      RECT 0.155 0.35 0.363 0.4 ;
      RECT 0.451 0.35 0.585 0.4 ;
      RECT 0.451 0.15 0.888 0.2 ;
      RECT 0.074 0.05 1.036 0.15 ;
    LAYER PO ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OAI33_0P5

MACRO SAEDRVT14_OA21_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.888 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.318 0.225 0.348 0.255 ;
      LAYER M2 ;
        RECT 0.241 0.223 0.397 0.257 ;
        RECT MASK 1 0.241 0.223 0.397 0.257 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.17 0.128 0.43 ;
        RECT 0.094 0.17 0.128 0.43 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.54 0.345 0.57 0.375 ;
      LAYER M2 ;
        RECT 0.463 0.343 0.619 0.377 ;
        RECT MASK 1 0.463 0.343 0.619 0.377 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.76 0.117 0.794 0.493 ;
        RECT MASK 1 0.76 0.117 0.794 0.493 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.93 0.647 ;
        RECT MASK 1 -0.042 0.553 0.93 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.93 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.93 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.39 0.454 0.72 0.488 ;
      RECT MASK 1 0.686 0.143 0.72 0.454 ;
      RECT MASK 1 0.612 0.109 0.72 0.143 ;
      RECT MASK 1 0.168 0.454 0.35 0.488 ;
      RECT MASK 1 0.316 0.414 0.35 0.454 ;
      RECT MASK 1 0.316 0.38 0.498 0.414 ;
      RECT MASK 1 0.538 0.237 0.572 0.414 ;
      RECT MASK 1 0.316 0.186 0.35 0.34 ;
      RECT MASK 1 0.168 0.112 0.572 0.146 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.962 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.814 0.55 ;
      RECT 0.074 0.4 0.296 0.45 ;
      RECT 0.666 0.4 0.814 0.45 ;
      RECT 0.296 0.2 0.444 0.25 ;
      RECT 0.074 0.05 0.444 0.2 ;
      RECT 0.666 0.15 0.814 0.2 ;
      RECT 0.518 0.05 0.814 0.15 ;
    LAYER PO ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OA21_U_0P5

MACRO SAEDRVT14_EO2_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.814 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.371 0.225 0.401 0.255 ;
      LAYER M2 ;
        RECT 0.345 0.223 0.601 0.257 ;
        RECT MASK 1 0.345 0.223 0.601 0.257 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.178 0.128 0.347 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.686 0.118 0.72 0.458 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.856 0.647 ;
        RECT MASK 1 -0.042 0.553 0.856 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.856 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.856 0.047 ;
    END
  END VSS
  OBS
    LAYER M2 ;
      RECT MASK 1 0.267 0.343 0.622 0.377 ;
    LAYER VIA1 ;
      RECT 0.548 0.345 0.578 0.375 ;
      RECT 0.293 0.345 0.323 0.375 ;
      RECT 0.449 0.285 0.479 0.315 ;
      RECT 0.209 0.285 0.239 0.315 ;
    LAYER M1 ;
      RECT MASK 1 0.228 0.45 0.66 0.488 ;
      RECT MASK 1 0.626 0.15 0.66 0.45 ;
      RECT MASK 1 0.312 0.112 0.66 0.15 ;
      RECT MASK 1 0.541 0.19 0.587 0.41 ;
      RECT MASK 1 0.15 0.361 0.241 0.395 ;
      RECT MASK 1 0.207 0.15 0.241 0.361 ;
      RECT MASK 1 0.15 0.112 0.241 0.15 ;
      RECT MASK 1 0.369 0.199 0.403 0.377 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.888 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.74 0.55 ;
      RECT 0.074 0.05 0.74 0.15 ;
    LAYER PO ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_EO2_0P5

MACRO SAEDRVT14_FDP_V2LP_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.702 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.152 0.128 0.443 ;
        RECT 0.094 0.152 0.128 0.443 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.354 0.285 1.384 0.315 ;
      LAYER M2 ;
        RECT 1.112 0.283 1.475 0.317 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.058 0.405 1.088 0.435 ;
      LAYER M2 ;
        RECT 0.961 0.403 1.185 0.437 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 1.5 0.091 1.534 0.507 ;
        RECT 1.5 0.091 1.534 0.507 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 0.553 1.744 0.647 ;
        RECT -0.042 0.553 1.744 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.046 1.744 0.048 ;
        RECT MASK 1 -0.042 -0.046 1.744 0.048 ;
    END
  END VSS
  OBS
    LAYER M2 ;
      RECT MASK 1 0.16 0.343 1.334 0.377 ;
      RECT MASK 1 0.294 0.223 1.266 0.257 ;
    LAYER VIA1 ;
      RECT 1.28 0.345 1.31 0.375 ;
      RECT 0.614 0.345 0.644 0.375 ;
      RECT 0.17 0.345 0.2 0.375 ;
      RECT 0.91 0.285 0.94 0.315 ;
      RECT 0.762 0.285 0.792 0.315 ;
      RECT 0.497 0.285 0.527 0.315 ;
      RECT 0.244 0.285 0.274 0.315 ;
      RECT 1.206 0.225 1.236 0.255 ;
      RECT 0.688 0.225 0.718 0.255 ;
      RECT 0.318 0.225 0.348 0.255 ;
      RECT 1.428 0.165 1.458 0.195 ;
      RECT 0.836 0.165 0.866 0.195 ;
    LAYER M1 ;
      RECT MASK 1 1.056 0.091 1.09 0.507 ;
      RECT MASK 1 0.316 0.41 0.35 0.507 ;
      RECT MASK 1 0.242 0.376 0.35 0.41 ;
      RECT MASK 1 0.242 0.091 0.276 0.376 ;
      RECT MASK 1 1.278 0.464 1.409 0.498 ;
      RECT MASK 1 1.278 0.137 1.312 0.464 ;
      RECT MASK 1 1.278 0.103 1.409 0.137 ;
      RECT MASK 1 0.67 0.464 0.868 0.498 ;
      RECT MASK 1 0.834 0.138 0.868 0.464 ;
      RECT MASK 1 0.59 0.104 0.868 0.138 ;
      RECT MASK 1 0.419 0.464 0.594 0.498 ;
      RECT MASK 1 0.419 0.222 0.453 0.464 ;
      RECT MASK 1 0.419 0.188 0.572 0.222 ;
      RECT MASK 1 1.204 0.123 1.238 0.477 ;
      RECT MASK 1 0.908 0.315 0.942 0.477 ;
      RECT MASK 1 0.908 0.281 1.013 0.315 ;
      RECT MASK 1 0.908 0.123 0.942 0.281 ;
      RECT MASK 1 0.168 0.233 0.202 0.477 ;
      RECT MASK 1 1.426 0.163 1.46 0.424 ;
      RECT MASK 1 1.352 0.256 1.386 0.424 ;
      RECT MASK 1 0.495 0.263 0.529 0.424 ;
      RECT MASK 1 0.612 0.206 0.646 0.422 ;
      RECT MASK 1 0.76 0.206 0.794 0.392 ;
      RECT MASK 1 0.686 0.206 0.72 0.392 ;
      RECT MASK 1 0.316 0.165 0.35 0.326 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.776 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 1.628 0.55 ;
      RECT 0.962 0.35 1.184 0.45 ;
      RECT 1.406 0.35 1.628 0.45 ;
      RECT 0.962 0.15 1.184 0.25 ;
      RECT 1.406 0.15 1.628 0.25 ;
      RECT 0.074 0.05 1.628 0.15 ;
    LAYER PO ;
      RECT 1.695 0 1.709 0.6 ;
      RECT 1.621 0 1.635 0.6 ;
      RECT 1.547 0 1.561 0.6 ;
      RECT 1.473 0 1.487 0.6 ;
      RECT 1.399 0 1.413 0.6 ;
      RECT 1.325 0 1.339 0.6 ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_FDP_V2LP_2

MACRO SAEDRVT14_FSDPQB_V2LP_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.924 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.327 0.345 0.357 0.375 ;
      LAYER M2 ;
        RECT 0.235 0.343 0.466 0.377 ;
        RECT MASK 1 0.235 0.343 0.466 0.377 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.429 0.285 0.459 0.315 ;
      LAYER M2 ;
        RECT 0.189 0.283 0.505 0.317 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.172 0.165 0.202 0.195 ;
        RECT 0.516 0.165 0.546 0.195 ;
      LAYER M2 ;
        RECT 0.151 0.163 0.555 0.197 ;
    END
  END SE
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.576 0.165 1.606 0.195 ;
      LAYER M2 ;
        RECT 1.554 0.163 1.79 0.197 ;
    END
  END CK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.722 0.102 1.756 0.488 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.966 0.647 ;
        RECT MASK 1 -0.042 0.553 1.966 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.966 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.966 0.047 ;
    END
  END VSS
  OBS
    LAYER M2 ;
      RECT MASK 1 0.76 0.343 1.564 0.377 ;
      RECT MASK 1 0.603 0.223 1.628 0.257 ;
    LAYER VIA1 ;
      RECT 1.433 0.345 1.463 0.375 ;
      RECT 1.021 0.345 1.051 0.375 ;
      RECT 0.765 0.345 0.795 0.375 ;
      RECT 1.653 0.285 1.683 0.315 ;
      RECT 1.284 0.285 1.314 0.315 ;
      RECT 0.922 0.285 0.952 0.315 ;
      RECT 0.679 0.285 0.709 0.315 ;
      RECT 1.502 0.225 1.532 0.255 ;
      RECT 1.117 0.225 1.147 0.255 ;
      RECT 0.605 0.225 0.635 0.255 ;
      RECT 1.359 0.165 1.389 0.195 ;
      RECT 1.21 0.165 1.24 0.195 ;
    LAYER M1 ;
      RECT MASK 1 0.288 0.458 0.569 0.498 ;
      RECT MASK 1 0.535 0.394 0.569 0.458 ;
      RECT MASK 1 0.612 0.395 0.646 0.488 ;
      RECT MASK 1 0.612 0.361 0.711 0.395 ;
      RECT MASK 1 0.677 0.102 0.711 0.361 ;
      RECT MASK 1 0.094 0.4 0.135 0.488 ;
      RECT MASK 1 0.094 0.366 0.28 0.4 ;
      RECT MASK 1 0.094 0.102 0.129 0.366 ;
      RECT MASK 1 0.246 0.263 0.28 0.366 ;
      RECT MASK 1 1.431 0.118 1.465 0.458 ;
      RECT MASK 1 1.357 0.118 1.391 0.458 ;
      RECT MASK 1 0.763 0.224 0.797 0.458 ;
      RECT MASK 1 1.014 0.263 1.06 0.425 ;
      RECT MASK 1 1.574 0.163 1.608 0.418 ;
      RECT MASK 1 0.915 0.263 0.961 0.418 ;
      RECT MASK 1 0.325 0.163 0.359 0.418 ;
      RECT MASK 1 1.651 0.175 1.685 0.4 ;
      RECT MASK 1 1.208 0.163 1.242 0.377 ;
      RECT MASK 1 1.115 0.199 1.149 0.377 ;
      RECT MASK 1 0.427 0.186 0.461 0.377 ;
      RECT MASK 1 0.169 0.163 0.204 0.326 ;
      RECT MASK 1 0.595 0.176 0.637 0.313 ;
      RECT MASK 1 0.509 0.163 0.555 0.313 ;
      RECT MASK 1 0.228 0.102 0.622 0.136 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.998 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 1.85 0.55 ;
      RECT 1.628 0.35 1.85 0.45 ;
      RECT 1.628 0.15 1.85 0.25 ;
      RECT 0.074 0.05 1.85 0.15 ;
    LAYER PO ;
      RECT 1.917 0 1.931 0.6 ;
      RECT 1.843 0 1.857 0.6 ;
      RECT 1.769 0 1.783 0.6 ;
      RECT 1.695 0 1.709 0.6 ;
      RECT 1.621 0 1.635 0.6 ;
      RECT 1.547 0 1.561 0.6 ;
      RECT 1.473 0 1.487 0.6 ;
      RECT 1.399 0 1.413 0.6 ;
      RECT 1.325 0 1.339 0.6 ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_FSDPQB_V2LP_2

MACRO SAEDRVT14_AO22_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.888 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.21 0.424 0.388 ;
        RECT 0.39 0.21 0.424 0.388 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.21 0.646 0.388 ;
        RECT MASK 1 0.612 0.21 0.646 0.388 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.235 0.276 0.389 ;
        RECT 0.242 0.235 0.276 0.389 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.111 0.128 0.388 ;
        RECT MASK 1 0.094 0.111 0.128 0.388 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.76 0.099 0.794 0.499 ;
        RECT MASK 1 0.76 0.099 0.794 0.499 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.93 0.647 ;
        RECT MASK 1 -0.042 0.553 0.93 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.93 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.93 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.094 0.442 0.683 0.476 ;
      RECT MASK 1 0.464 0.354 0.572 0.388 ;
      RECT MASK 1 0.686 0.165 0.72 0.363 ;
      RECT MASK 1 0.538 0.165 0.572 0.354 ;
      RECT MASK 1 0.302 0.127 0.72 0.165 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.962 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.814 0.55 ;
      RECT 0.074 0.4 0.37 0.45 ;
      RECT 0.074 0.35 0.222 0.4 ;
      RECT 0.074 0.15 0.37 0.25 ;
      RECT 0.074 0.05 0.814 0.15 ;
    LAYER PO ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AO22_0P5

MACRO SAEDRVT14_OA221_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.814 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.209 0.276 0.418 ;
        RECT 0.242 0.209 0.276 0.418 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.115 0.405 0.145 0.435 ;
      LAYER M2 ;
        RECT -0.007 0.403 0.229 0.437 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.245 0.35 0.393 ;
        RECT MASK 1 0.316 0.245 0.35 0.393 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 0.263 0.424 0.418 ;
        RECT MASK 1 0.39 0.263 0.424 0.418 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.526 0.285 0.556 0.315 ;
      LAYER M2 ;
        RECT 0.437 0.283 0.673 0.317 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.686 0.114 0.72 0.496 ;
        RECT MASK 1 0.686 0.114 0.72 0.496 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.856 0.647 ;
        RECT MASK 1 -0.042 0.553 0.856 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.856 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.856 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.228 0.458 0.64 0.496 ;
      RECT MASK 1 0.606 0.14 0.64 0.458 ;
      RECT MASK 1 0.533 0.102 0.64 0.14 ;
      RECT MASK 1 0.107 0.288 0.153 0.488 ;
      RECT MASK 1 0.519 0.254 0.565 0.377 ;
      RECT MASK 1 0.304 0.18 0.544 0.214 ;
      RECT MASK 1 0.085 0.14 0.123 0.207 ;
      RECT MASK 1 0.085 0.102 0.46 0.14 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.888 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.74 0.55 ;
      RECT 0.074 0.15 0.592 0.2 ;
      RECT 0.074 0.05 0.74 0.15 ;
    LAYER PO ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OA221_U_0P5

MACRO SAEDRVT14_AO31_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.036 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.542 0.225 0.572 0.255 ;
      LAYER M2 ;
        RECT 0.405 0.223 0.619 0.257 ;
        RECT MASK 1 0.405 0.223 0.619 0.257 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.26 0.35 0.414 ;
        RECT MASK 1 0.316 0.26 0.35 0.414 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.162 0.128 0.457 ;
        RECT MASK 1 0.094 0.162 0.128 0.457 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.688 0.225 0.718 0.255 ;
      LAYER M2 ;
        RECT 0.678 0.223 0.908 0.257 ;
        RECT MASK 1 0.678 0.223 0.908 0.257 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.908 0.095 0.942 0.507 ;
        RECT MASK 1 0.908 0.095 0.942 0.507 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.078 0.647 ;
        RECT MASK 1 -0.042 0.553 1.078 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.078 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.078 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.168 0.454 0.72 0.488 ;
      RECT MASK 1 0.76 0.451 0.868 0.485 ;
      RECT MASK 1 0.834 0.145 0.868 0.451 ;
      RECT MASK 1 0.612 0.111 0.868 0.145 ;
      RECT MASK 1 0.686 0.214 0.72 0.414 ;
      RECT MASK 1 0.54 0.217 0.574 0.414 ;
      RECT MASK 1 0.316 0.179 0.498 0.213 ;
      RECT MASK 1 0.316 0.153 0.35 0.179 ;
      RECT MASK 1 0.168 0.105 0.35 0.153 ;
      RECT MASK 1 0.39 0.105 0.572 0.139 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.11 0.6 ;
    LAYER DIFF ;
      RECT 0.518 0.4 0.962 0.55 ;
      RECT 0.666 0.35 0.962 0.4 ;
      RECT 0.074 0.4 0.444 0.55 ;
      RECT 0.296 0.35 0.444 0.4 ;
      RECT 0.518 0.2 0.666 0.25 ;
      RECT 0.074 0.15 0.666 0.2 ;
      RECT 0.814 0.15 0.962 0.2 ;
      RECT 0.074 0.05 0.962 0.15 ;
    LAYER PO ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AO31_1

MACRO SAEDRVT14_FDPSYNSBQ_V2_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.072 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.316 0.169 0.35 0.435 ;
        RECT 0.316 0.169 0.35 0.435 ;
    END
  END D
  PIN SD
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.206 0.202 0.392 ;
        RECT 0.168 0.206 0.202 0.392 ;
    END
  END SD
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.354 0.165 1.384 0.195 ;
      LAYER M2 ;
        RECT 1.337 0.163 1.623 0.197 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.876 0.225 1.906 0.255 ;
      LAYER M2 ;
        RECT 1.72 0.223 2.154 0.257 ;
        RECT MASK 1 1.72 0.223 2.154 0.257 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 2.114 0.647 ;
        RECT MASK 1 -0.042 0.553 2.114 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.048 2.114 0.047 ;
        RECT MASK 1 -0.042 -0.048 2.114 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 1.5 0.123 1.534 0.477 ;
      RECT MASK 1 1.204 0.163 1.238 0.477 ;
      RECT MASK 1 0.612 0.233 0.646 0.477 ;
      RECT MASK 1 1.648 0.163 1.682 0.435 ;
      RECT MASK 1 1.352 0.163 1.386 0.435 ;
      RECT MASK 1 0.77 0.269 0.804 0.43 ;
      RECT MASK 1 0.858 0.268 0.892 0.429 ;
      RECT MASK 1 1.056 0.17 1.09 0.392 ;
      RECT MASK 1 0.464 0.169 0.498 0.326 ;
    LAYER M2 ;
      RECT MASK 1 0.576 0.343 1.55 0.377 ;
      RECT MASK 1 0.442 0.223 1.482 0.257 ;
    LAYER VIA1 ;
      RECT 1.502 0.345 1.532 0.375 ;
      RECT 0.86 0.345 0.89 0.375 ;
      RECT 0.614 0.345 0.644 0.375 ;
      RECT 1.65 0.285 1.68 0.315 ;
      RECT 1.206 0.285 1.236 0.315 ;
      RECT 1.058 0.285 1.088 0.315 ;
      RECT 0.772 0.285 0.802 0.315 ;
      RECT 0.54 0.285 0.57 0.315 ;
      RECT 1.428 0.225 1.458 0.255 ;
      RECT 0.952 0.225 0.982 0.255 ;
      RECT 0.466 0.225 0.496 0.255 ;
    LAYER NWELL ;
      RECT -0.074 0.3 2.146 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 1.998 0.55 ;
      RECT 1.48 0.4 1.998 0.45 ;
      RECT 1.628 0.35 1.998 0.4 ;
      RECT 1.628 0.2 1.998 0.25 ;
      RECT 1.332 0.15 1.998 0.2 ;
      RECT 0.444 0.05 1.998 0.15 ;
      RECT 0.074 0.05 0.37 0.15 ;
    LAYER PO ;
      RECT 2.065 0 2.079 0.6 ;
      RECT 1.991 0 2.005 0.6 ;
      RECT 1.917 0 1.931 0.6 ;
      RECT 1.843 0 1.857 0.6 ;
      RECT 1.769 0 1.783 0.6 ;
      RECT 1.695 0 1.709 0.6 ;
      RECT 1.621 0 1.635 0.6 ;
      RECT 1.547 0 1.561 0.6 ;
      RECT 1.473 0 1.487 0.6 ;
      RECT 1.399 0 1.413 0.6 ;
      RECT 1.325 0 1.339 0.6 ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_FDPSYNSBQ_V2_4

MACRO SAEDRVT14_LDNQ_V1_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.11 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.092 0.202 0.503 ;
        RECT 0.168 0.092 0.202 0.503 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.762 0.165 0.792 0.195 ;
      LAYER M2 ;
        RECT 0.456 0.163 0.794 0.197 ;
    END
  END G
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.982 0.102 1.016 0.497 ;
        RECT MASK 1 0.982 0.102 1.016 0.497 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.152 0.647 ;
        RECT MASK 1 -0.042 0.553 1.152 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.152 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.152 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.612 0.118 0.646 0.458 ;
      RECT MASK 1 0.478 0.156 0.512 0.419 ;
      RECT MASK 1 0.332 0.283 0.376 0.416 ;
      RECT MASK 1 0.908 0.102 0.942 0.363 ;
      RECT MASK 1 0.76 0.118 0.794 0.287 ;
    LAYER M2 ;
      RECT MASK 1 0.449 0.343 0.694 0.377 ;
      RECT MASK 1 0.398 0.223 0.791 0.257 ;
      RECT MASK 1 0.303 0.103 0.967 0.137 ;
    LAYER VIA1 ;
      RECT 0.614 0.345 0.644 0.375 ;
      RECT 0.48 0.345 0.51 0.375 ;
      RECT 0.836 0.285 0.866 0.315 ;
      RECT 0.344 0.285 0.374 0.315 ;
      RECT 0.688 0.225 0.718 0.255 ;
      RECT 0.413 0.225 0.443 0.255 ;
      RECT 0.91 0.105 0.94 0.135 ;
      RECT 0.547 0.105 0.577 0.135 ;
      RECT 0.318 0.105 0.348 0.135 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.184 0.6 ;
    LAYER DIFF ;
      RECT 0.296 0.45 1.036 0.55 ;
      RECT 0.888 0.35 1.036 0.45 ;
      RECT 0.074 0.35 0.222 0.55 ;
      RECT 0.074 0.15 0.222 0.25 ;
      RECT 0.888 0.15 1.036 0.25 ;
      RECT 0.074 0.05 1.036 0.15 ;
    LAYER PO ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_LDNQ_V1_1

MACRO SAEDRVT14_OAI311_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.962 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.234 0.35 0.418 ;
        RECT MASK 1 0.316 0.234 0.35 0.418 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.237 0.276 0.513 ;
        RECT MASK 1 0.242 0.237 0.276 0.513 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.24 0.128 0.458 ;
        RECT MASK 1 0.094 0.24 0.128 0.458 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.464 0.2 0.498 0.377 ;
        RECT MASK 1 0.464 0.2 0.498 0.377 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.222 0.424 0.397 ;
        RECT 0.39 0.222 0.424 0.397 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.834 0.107 0.868 0.496 ;
        RECT 0.834 0.107 0.868 0.496 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.004 0.647 ;
        RECT MASK 1 -0.042 0.553 1.004 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.004 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.004 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.684 0.319 0.722 0.496 ;
      RECT MASK 1 0.684 0.285 0.792 0.319 ;
      RECT MASK 1 0.684 0.107 0.722 0.285 ;
      RECT MASK 1 0.367 0.458 0.574 0.496 ;
      RECT MASK 1 0.536 0.319 0.574 0.458 ;
      RECT MASK 1 0.536 0.285 0.644 0.319 ;
      RECT MASK 1 0.536 0.107 0.574 0.285 ;
      RECT MASK 1 0.15 0.102 0.388 0.14 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.036 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.888 0.55 ;
      RECT 0.155 0.4 0.303 0.45 ;
      RECT 0.229 0.35 0.303 0.4 ;
      RECT 0.451 0.15 0.525 0.2 ;
      RECT 0.074 0.05 0.888 0.15 ;
    LAYER PO ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OAI311_0P5

MACRO SAEDRVT14_TIE0_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.814 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.686 0.112 0.72 0.488 ;
        RECT MASK 1 0.337 0.45 0.72 0.488 ;
        RECT MASK 1 0.337 0.369 0.375 0.45 ;
        RECT MASK 1 0.686 0.15 0.72 0.45 ;
        RECT MASK 1 0.315 0.15 0.353 0.207 ;
        RECT MASK 1 0.315 0.112 0.72 0.15 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.856 0.647 ;
        RECT MASK 1 -0.042 0.553 0.856 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.856 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.856 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.15 0.422 0.281 0.46 ;
      RECT MASK 1 0.247 0.311 0.281 0.422 ;
      RECT MASK 1 0.247 0.265 0.371 0.311 ;
      RECT MASK 1 0.129 0.15 0.175 0.329 ;
      RECT MASK 1 0.129 0.112 0.232 0.15 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.888 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.74 0.55 ;
      RECT 0.074 0.35 0.222 0.4 ;
      RECT 0.074 0.2 0.222 0.25 ;
      RECT 0.074 0.05 0.74 0.2 ;
    LAYER PO ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_TIE0_4

MACRO SAEDRVT14_TIE1_V1_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.37 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.173 0.276 0.475 ;
        RECT MASK 1 0.15 0.437 0.276 0.475 ;
        RECT MASK 1 0.242 0.173 0.276 0.437 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.412 0.647 ;
        RECT MASK 1 -0.042 0.553 0.412 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.412 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.412 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.129 0.15 0.175 0.361 ;
      RECT MASK 1 0.129 0.112 0.213 0.15 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.444 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.296 0.55 ;
      RECT 0.074 0.05 0.296 0.2 ;
    LAYER PO ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_TIE1_V1_2

MACRO SAEDRVT14_EO3_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.702 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.762 0.345 0.792 0.375 ;
      LAYER M2 ;
        RECT MASK 1 0.748 0.343 1.146 0.377 ;
        RECT 0.748 0.343 1.146 0.377 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.344 0.225 0.374 0.255 ;
      LAYER M2 ;
        RECT 0.304 0.223 0.679 0.257 ;
        RECT MASK 1 0.304 0.223 0.679 0.257 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.181 0.128 0.405 ;
        RECT 0.094 0.181 0.128 0.405 ;
    END
  END A3
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.574 0.118 1.608 0.458 ;
        RECT MASK 1 1.574 0.118 1.608 0.458 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.744 0.647 ;
        RECT MASK 1 -0.042 0.553 1.744 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.744 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.744 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.834 0.165 0.868 0.505 ;
      RECT MASK 1 0.95 0.458 1.236 0.496 ;
      RECT MASK 1 1.202 0.136 1.236 0.458 ;
      RECT MASK 1 0.905 0.102 1.236 0.136 ;
      RECT MASK 1 0.241 0.458 0.646 0.496 ;
      RECT MASK 1 0.612 0.14 0.646 0.458 ;
      RECT MASK 1 0.282 0.102 0.646 0.14 ;
      RECT MASK 1 1.426 0.318 1.46 0.458 ;
      RECT MASK 1 1.426 0.284 1.534 0.318 ;
      RECT MASK 1 1.426 0.118 1.46 0.284 ;
      RECT MASK 1 1.278 0.318 1.312 0.458 ;
      RECT MASK 1 1.278 0.284 1.386 0.318 ;
      RECT MASK 1 1.278 0.118 1.312 0.284 ;
      RECT MASK 1 0.76 0.263 0.794 0.437 ;
      RECT MASK 1 0.922 0.163 0.956 0.418 ;
      RECT MASK 1 0.686 0.158 0.72 0.418 ;
      RECT MASK 1 0.538 0.18 0.572 0.418 ;
      RECT MASK 1 0.416 0.199 0.45 0.418 ;
      RECT MASK 1 0.268 0.185 0.302 0.418 ;
      RECT MASK 1 0.168 0.361 0.212 0.395 ;
      RECT MASK 1 0.178 0.141 0.212 0.361 ;
      RECT MASK 1 0.121 0.103 0.212 0.141 ;
      RECT MASK 1 1.075 0.177 1.109 0.377 ;
      RECT MASK 1 0.996 0.199 1.03 0.377 ;
      RECT MASK 1 0.342 0.199 0.376 0.377 ;
    LAYER M2 ;
      RECT MASK 1 0.248 0.343 0.589 0.377 ;
      RECT MASK 1 0.813 0.223 1.207 0.257 ;
    LAYER VIA1 ;
      RECT 0.54 0.345 0.57 0.375 ;
      RECT 0.27 0.345 0.3 0.375 ;
      RECT 0.998 0.285 1.028 0.315 ;
      RECT 0.614 0.285 0.644 0.315 ;
      RECT 0.418 0.285 0.448 0.315 ;
      RECT 0.18 0.285 0.21 0.315 ;
      RECT 1.077 0.225 1.107 0.255 ;
      RECT 0.836 0.225 0.866 0.255 ;
      RECT 0.924 0.165 0.954 0.195 ;
      RECT 0.688 0.165 0.718 0.195 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.776 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 1.628 0.55 ;
      RECT 1.399 0.4 1.473 0.45 ;
      RECT 0.363 0.15 0.437 0.2 ;
      RECT 0.511 0.15 0.599 0.2 ;
      RECT 1.399 0.15 1.473 0.2 ;
      RECT 0.074 0.05 1.628 0.15 ;
    LAYER PO ;
      RECT 1.695 0 1.709 0.6 ;
      RECT 1.621 0 1.635 0.6 ;
      RECT 1.547 0 1.561 0.6 ;
      RECT 1.473 0 1.487 0.6 ;
      RECT 1.399 0 1.413 0.6 ;
      RECT 1.325 0 1.339 0.6 ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_EO3_0P5

MACRO SAEDRVT14_OAI311_0P75
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.962 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.316 0.234 0.35 0.418 ;
        RECT MASK 1 0.316 0.234 0.35 0.418 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.237 0.276 0.505 ;
        RECT 0.242 0.237 0.276 0.505 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.24 0.128 0.458 ;
        RECT MASK 1 0.094 0.24 0.128 0.458 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.464 0.2 0.498 0.377 ;
        RECT 0.464 0.2 0.498 0.377 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 0.222 0.424 0.397 ;
        RECT MASK 1 0.39 0.222 0.424 0.397 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.834 0.107 0.868 0.496 ;
        RECT 0.834 0.107 0.868 0.496 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.004 0.647 ;
        RECT MASK 1 -0.042 0.553 1.004 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.004 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.004 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.684 0.319 0.722 0.496 ;
      RECT MASK 1 0.684 0.285 0.792 0.319 ;
      RECT MASK 1 0.684 0.107 0.722 0.285 ;
      RECT MASK 1 0.367 0.458 0.574 0.496 ;
      RECT MASK 1 0.536 0.319 0.574 0.458 ;
      RECT MASK 1 0.536 0.285 0.644 0.319 ;
      RECT MASK 1 0.536 0.107 0.574 0.285 ;
      RECT MASK 1 0.15 0.102 0.388 0.14 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.036 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.888 0.55 ;
      RECT 0.155 0.4 0.303 0.45 ;
      RECT 0.229 0.35 0.303 0.4 ;
      RECT 0.451 0.15 0.525 0.2 ;
      RECT 0.074 0.05 0.888 0.15 ;
    LAYER PO ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OAI311_0P75

MACRO SAEDRVT14_EO2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.814 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.371 0.225 0.401 0.255 ;
      LAYER M2 ;
        RECT 0.345 0.223 0.601 0.257 ;
        RECT MASK 1 0.345 0.223 0.601 0.257 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.088 0.175 0.122 0.334 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.686 0.118 0.72 0.458 ;
        RECT 0.686 0.118 0.72 0.458 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.856 0.647 ;
        RECT MASK 1 -0.042 0.553 0.856 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.856 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.856 0.047 ;
    END
  END VSS
  OBS
    LAYER M2 ;
      RECT MASK 1 0.267 0.343 0.622 0.377 ;
    LAYER VIA1 ;
      RECT 0.548 0.345 0.578 0.375 ;
      RECT 0.293 0.345 0.323 0.375 ;
      RECT 0.449 0.285 0.479 0.315 ;
      RECT 0.209 0.285 0.239 0.315 ;
    LAYER M1 ;
      RECT MASK 1 0.541 0.19 0.587 0.41 ;
      RECT MASK 1 0.15 0.361 0.241 0.395 ;
      RECT MASK 1 0.207 0.15 0.241 0.361 ;
      RECT MASK 1 0.15 0.112 0.241 0.15 ;
      RECT MASK 1 0.369 0.199 0.403 0.377 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.888 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.74 0.55 ;
      RECT 0.592 0.35 0.74 0.45 ;
      RECT 0.592 0.15 0.74 0.25 ;
      RECT 0.074 0.05 0.74 0.15 ;
    LAYER PO ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_EO2_1

MACRO SAEDRVT14_ND2_MM_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.518 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.316 0.264 0.35 0.477 ;
        RECT 0.316 0.264 0.35 0.477 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.182 0.202 0.437 ;
        RECT 0.168 0.182 0.202 0.437 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.176 0.276 0.509 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.56 0.647 ;
        RECT MASK 1 -0.042 0.553 0.56 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.56 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.56 0.047 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.3 0.592 0.6 ;
    LAYER DIFF ;
      RECT 0.148 0.45 0.37 0.55 ;
      RECT 0.074 0.05 0.444 0.15 ;
    LAYER PO ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_ND2_MM_0P5

MACRO SAEDRVT14_AO222_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.332 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.908 0.19 0.942 0.344 ;
        RECT 0.908 0.19 0.942 0.344 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 1.058 0.285 1.088 0.315 ;
      LAYER M2 ;
        RECT 0.99 0.283 1.141 0.317 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.76 0.19 0.794 0.344 ;
        RECT 0.76 0.19 0.794 0.344 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.54 0.345 0.57 0.375 ;
      LAYER M2 ;
        RECT 0.481 0.343 0.631 0.377 ;
        RECT MASK 1 0.481 0.343 0.631 0.377 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.316 0.27 0.35 0.424 ;
        RECT 0.316 0.27 0.35 0.424 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.104 0.128 0.474 ;
        RECT MASK 1 0.094 0.104 0.128 0.474 ;
    END
  END C2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.204 0.117 1.238 0.493 ;
        RECT MASK 1 1.204 0.117 1.238 0.493 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.374 0.647 ;
        RECT MASK 1 -0.042 0.553 1.374 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.374 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.374 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.168 0.464 0.72 0.498 ;
      RECT MASK 1 0.76 0.461 1.016 0.495 ;
      RECT MASK 1 0.76 0.421 0.794 0.461 ;
      RECT MASK 1 0.612 0.387 0.794 0.421 ;
      RECT MASK 1 0.538 0.176 0.572 0.421 ;
      RECT MASK 1 0.834 0.384 1.164 0.418 ;
      RECT MASK 1 0.834 0.15 0.868 0.384 ;
      RECT MASK 1 1.13 0.117 1.164 0.384 ;
      RECT MASK 1 0.39 0.116 0.868 0.15 ;
      RECT MASK 1 1.056 0.19 1.09 0.344 ;
      RECT MASK 1 0.612 0.21 0.72 0.258 ;
      RECT MASK 1 0.316 0.19 0.498 0.224 ;
      RECT MASK 1 0.316 0.146 0.35 0.19 ;
      RECT MASK 1 0.168 0.112 0.35 0.146 ;
      RECT MASK 1 0.908 0.116 1.063 0.15 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.406 0.6 ;
    LAYER DIFF ;
      RECT 0.518 0.45 1.258 0.55 ;
      RECT 0.518 0.4 0.814 0.45 ;
      RECT 1.11 0.4 1.258 0.45 ;
      RECT 0.518 0.35 0.666 0.4 ;
      RECT 0.074 0.4 0.444 0.55 ;
      RECT 0.296 0.35 0.444 0.4 ;
      RECT 0.666 0.2 0.814 0.25 ;
      RECT 0.296 0.15 0.814 0.2 ;
      RECT 1.11 0.15 1.258 0.2 ;
      RECT 0.296 0.05 1.258 0.15 ;
      RECT 0.074 0.05 0.222 0.25 ;
    LAYER PO ;
      RECT 1.325 0 1.339 0.6 ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AO222_U_0P5

MACRO SAEDRVT14_AN2_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.666 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.18 0.276 0.418 ;
        RECT MASK 1 0.242 0.18 0.276 0.418 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.18 0.128 0.418 ;
        RECT MASK 1 0.094 0.18 0.128 0.418 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.443 0.424 0.477 ;
        RECT MASK 1 0.39 0.409 0.573 0.443 ;
        RECT MASK 1 0.39 0.123 0.424 0.409 ;
        RECT 0.39 0.123 0.424 0.477 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.708 0.647 ;
        RECT MASK 1 -0.042 0.553 0.708 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.708 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.708 0.047 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.3 0.74 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.592 0.55 ;
      RECT 0.074 0.05 0.518 0.15 ;
    LAYER PO ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AN2_0P5

MACRO SAEDRVT14_MUXI2_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.888 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.168 0.123 0.202 0.326 ;
        RECT 0.168 0.123 0.202 0.326 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.464 0.176 0.498 0.424 ;
        RECT 0.464 0.176 0.498 0.424 ;
    END
  END D1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 0.176 0.424 0.424 ;
        RECT MASK 1 0.39 0.176 0.424 0.424 ;
    END
  END S
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.76 0.123 0.794 0.477 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.046 0.553 0.93 0.647 ;
        RECT MASK 1 -0.046 0.553 0.93 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.046 -0.047 0.93 0.047 ;
        RECT MASK 1 -0.046 -0.047 0.93 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.612 0.318 0.646 0.477 ;
      RECT MASK 1 0.612 0.279 0.695 0.318 ;
      RECT MASK 1 0.612 0.123 0.646 0.279 ;
    LAYER NWELL ;
      RECT -0.078 0.3 0.962 0.6 ;
    LAYER DIFF ;
      RECT 0.07 0.45 0.814 0.55 ;
      RECT 0.07 0.05 0.814 0.15 ;
    LAYER PO ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_MUXI2_0P5

MACRO SAEDRVT14_OA21B_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.888 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.204 0.225 0.234 0.255 ;
      LAYER M2 ;
        RECT 0.159 0.223 0.314 0.257 ;
        RECT MASK 1 0.159 0.223 0.314 0.257 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.199 0.128 0.442 ;
        RECT MASK 1 0.094 0.199 0.128 0.442 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.466 0.165 0.496 0.195 ;
      LAYER M2 ;
        RECT 0.455 0.163 0.626 0.197 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.76 0.085 0.794 0.459 ;
        RECT 0.76 0.085 0.794 0.459 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 0.553 0.93 0.647 ;
        RECT -0.042 0.553 0.93 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.93 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.93 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.594 0.443 0.697 0.488 ;
      RECT MASK 1 0.651 0.15 0.697 0.443 ;
      RECT MASK 1 0.594 0.112 0.697 0.15 ;
      RECT MASK 1 0.459 0.396 0.499 0.488 ;
      RECT MASK 1 0.459 0.395 0.591 0.396 ;
      RECT MASK 1 0.399 0.361 0.591 0.395 ;
      RECT MASK 1 0.399 0.088 0.433 0.361 ;
      RECT MASK 1 0.499 0.36 0.591 0.361 ;
      RECT MASK 1 0.557 0.192 0.591 0.36 ;
      RECT MASK 1 0.216 0.447 0.359 0.485 ;
      RECT MASK 1 0.325 0.154 0.359 0.447 ;
      RECT MASK 1 0.138 0.112 0.359 0.154 ;
      RECT MASK 1 0.195 0.199 0.241 0.352 ;
      RECT MASK 1 0.464 0.148 0.498 0.313 ;
      RECT 0.464 0.148 0.498 0.313 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.962 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.814 0.55 ;
      RECT 0.518 0.15 0.666 0.2 ;
      RECT 0.074 0.05 0.814 0.15 ;
    LAYER PO ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_OA21B_U_0P5

MACRO SAEDRVT14_NR2B_U_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.814 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.18 0.128 0.331 ;
        RECT MASK 1 0.094 0.18 0.128 0.331 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 0.142 0.424 0.329 ;
        RECT MASK 1 0.39 0.142 0.424 0.329 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.686 0.091 0.72 0.459 ;
        RECT MASK 1 0.686 0.091 0.72 0.459 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 0.553 0.856 0.647 ;
        RECT -0.042 0.553 0.856 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.856 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.856 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.52 0.443 0.623 0.488 ;
      RECT MASK 1 0.577 0.15 0.623 0.443 ;
      RECT MASK 1 0.52 0.112 0.623 0.15 ;
      RECT MASK 1 0.242 0.453 0.361 0.487 ;
      RECT MASK 1 0.316 0.398 0.35 0.453 ;
      RECT MASK 1 0.316 0.364 0.517 0.398 ;
      RECT MASK 1 0.316 0.114 0.35 0.364 ;
      RECT MASK 1 0.483 0.192 0.517 0.364 ;
      RECT MASK 1 0.168 0.392 0.202 0.426 ;
      RECT MASK 1 0.138 0.358 0.276 0.392 ;
      RECT MASK 1 0.242 0.15 0.276 0.358 ;
      RECT MASK 1 0.14 0.112 0.276 0.15 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.888 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.74 0.55 ;
      RECT 0.074 0.05 0.74 0.15 ;
    LAYER PO ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_NR2B_U_0P5

MACRO SAEDRVT14_NR2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.37 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.1 0.276 0.337 ;
        RECT 0.242 0.1 0.276 0.337 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.159 0.128 0.445 ;
        RECT 0.094 0.159 0.128 0.445 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.425 0.276 0.469 ;
        RECT MASK 1 0.168 0.391 0.276 0.425 ;
        RECT MASK 1 0.168 0.089 0.202 0.391 ;
        RECT 0.168 0.089 0.202 0.425 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 0.553 0.392 0.647 ;
        RECT -0.042 0.553 0.392 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT MASK 1 -0.042 -0.047 0.392 0.047 ;
        RECT -0.042 -0.047 0.392 0.047 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.299 0.424 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.296 0.55 ;
      RECT 0.074 0.05 0.296 0.15 ;
    LAYER PO ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_NR2_1

MACRO SAEDRVT14_ND3B_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.888 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.134 0.285 0.164 0.315 ;
      LAYER M2 ;
        RECT -0.026 0.283 0.176 0.317 ;
    END
  END A
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.339 0.345 0.369 0.375 ;
      LAYER M2 ;
        RECT MASK 1 0.169 0.343 0.371 0.377 ;
        RECT 0.169 0.343 0.371 0.377 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.41 0.285 0.44 0.315 ;
      LAYER M2 ;
        RECT 0.407 0.283 0.609 0.317 ;
    END
  END B2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.76 0.119 0.794 0.459 ;
        RECT MASK 1 0.76 0.119 0.794 0.459 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.93 0.647 ;
        RECT MASK 1 -0.042 0.553 0.93 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.93 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.93 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.596 0.45 0.699 0.488 ;
      RECT MASK 1 0.653 0.15 0.699 0.45 ;
      RECT MASK 1 0.612 0.112 0.699 0.15 ;
      RECT MASK 1 0.408 0.2 0.442 0.423 ;
      RECT MASK 1 0.148 0.389 0.3 0.423 ;
      RECT MASK 1 0.266 0.204 0.3 0.389 ;
      RECT MASK 1 0.148 0.17 0.3 0.204 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.962 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.814 0.55 ;
      RECT 0.074 0.4 0.222 0.45 ;
      RECT 0.518 0.35 0.666 0.45 ;
      RECT 0.074 0.15 0.363 0.2 ;
      RECT 0.074 0.05 0.814 0.15 ;
    LAYER PO ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_ND3B_0P5

MACRO SAEDRVT14_ND3_ECO_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.258 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.202 0.276 0.374 ;
        RECT 0.242 0.202 0.276 0.374 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.373 0.345 0.403 0.375 ;
      LAYER M2 ;
        RECT 0.254 0.343 0.506 0.377 ;
        RECT MASK 1 0.254 0.343 0.506 0.377 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.594 0.345 0.624 0.375 ;
      LAYER M2 ;
        RECT 0.592 0.343 0.85 0.377 ;
        RECT MASK 1 0.592 0.343 0.85 0.377 ;
    END
  END A3
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.834 0.102 0.868 0.498 ;
        RECT MASK 1 0.834 0.464 0.932 0.498 ;
        RECT MASK 1 0.834 0.152 0.868 0.464 ;
        RECT MASK 1 0.834 0.102 0.932 0.152 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.3 0.647 ;
        RECT MASK 1 -0.042 0.553 1.3 0.647 ;
        RECT MASK 1 0.094 0.414 0.128 0.553 ;
        RECT MASK 1 0.464 0.414 0.498 0.553 ;
        RECT MASK 1 0.686 0.451 0.72 0.553 ;
        RECT MASK 1 1.056 0.451 1.09 0.553 ;
        RECT MASK 1 0.686 0.414 0.794 0.451 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.3 0.047 ;
        RECT MASK 1 0.686 0.123 0.794 0.16 ;
        RECT MASK 1 1.056 0.047 1.09 0.165 ;
        RECT MASK 1 0.686 0.047 0.72 0.123 ;
        RECT MASK 1 -0.042 -0.047 1.3 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 1.13 0.092 1.164 0.511 ;
      RECT MASK 1 0.538 0.448 0.646 0.498 ;
      RECT MASK 1 0.168 0.463 0.389 0.497 ;
      RECT MASK 1 0.168 0.261 0.202 0.463 ;
      RECT MASK 1 0.094 0.227 0.202 0.261 ;
      RECT MASK 1 0.094 0.088 0.128 0.227 ;
      RECT MASK 1 0.982 0.088 1.016 0.488 ;
      RECT MASK 1 0.371 0.202 0.405 0.391 ;
      RECT MASK 1 0.592 0.202 0.626 0.382 ;
      RECT MASK 1 0.908 0.202 0.942 0.374 ;
      RECT MASK 1 0.464 0.136 0.498 0.207 ;
      RECT MASK 1 0.464 0.102 0.594 0.136 ;
      RECT MASK 1 0.168 0.102 0.35 0.136 ;
    LAYER M2 ;
      RECT MASK 1 0.159 0.463 1.171 0.497 ;
    LAYER VIA1 ;
      RECT 1.132 0.465 1.162 0.495 ;
      RECT 0.583 0.465 0.613 0.495 ;
      RECT 0.339 0.465 0.369 0.495 ;
      RECT 0.195 0.465 0.225 0.495 ;
      RECT 0.984 0.285 1.014 0.315 ;
      RECT 0.91 0.285 0.94 0.315 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.332 0.6 ;
    LAYER DIFF ;
      RECT 0.962 0.35 1.11 0.55 ;
      RECT 0.74 0.35 0.888 0.55 ;
      RECT 0.518 0.35 0.666 0.55 ;
      RECT 0.296 0.35 0.444 0.55 ;
      RECT 0.074 0.4 0.222 0.55 ;
      RECT 0.74 0.05 0.888 0.25 ;
      RECT 0.296 0.05 0.444 0.25 ;
      RECT 0.074 0.05 0.222 0.25 ;
      RECT 0.518 0.05 0.666 0.2 ;
      RECT 0.962 0.05 1.11 0.15 ;
    LAYER PO ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_ND3_ECO_1

MACRO SAEDRVT14_AOI31_0P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.814 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.205 0.276 0.418 ;
        RECT 0.242 0.205 0.276 0.418 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.17 0.105 0.2 0.135 ;
      LAYER M2 ;
        RECT MASK 1 0.082 0.103 0.352 0.137 ;
        RECT 0.082 0.103 0.352 0.137 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.096 0.405 0.126 0.435 ;
      LAYER M2 ;
        RECT -0.032 0.403 0.204 0.437 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.316 0.199 0.35 0.391 ;
        RECT 0.316 0.199 0.35 0.391 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.686 0.119 0.72 0.459 ;
        RECT 0.686 0.119 0.72 0.459 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.856 0.647 ;
        RECT MASK 1 -0.042 0.553 0.856 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.856 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.856 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.15 0.458 0.35 0.496 ;
      RECT MASK 1 0.52 0.443 0.623 0.488 ;
      RECT MASK 1 0.577 0.15 0.623 0.443 ;
      RECT MASK 1 0.52 0.112 0.623 0.15 ;
      RECT MASK 1 0.094 0.158 0.128 0.444 ;
      RECT MASK 1 0.39 0.358 0.517 0.392 ;
      RECT MASK 1 0.483 0.192 0.517 0.358 ;
      RECT MASK 1 0.39 0.154 0.424 0.358 ;
      RECT MASK 1 0.312 0.116 0.424 0.154 ;
      RECT MASK 1 0.168 0.088 0.202 0.377 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.888 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.74 0.55 ;
      RECT 0.363 0.35 0.444 0.45 ;
      RECT 0.289 0.2 0.363 0.25 ;
      RECT 0.155 0.15 0.363 0.2 ;
      RECT 0.074 0.05 0.74 0.15 ;
    LAYER PO ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AOI31_0P5

MACRO SAEDRVT14_ND2B_0P75
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.036 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.144 0.128 0.466 ;
        RECT 0.094 0.144 0.128 0.466 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.39 0.193 0.424 0.414 ;
        RECT MASK 1 0.39 0.193 0.424 0.414 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.836 0.225 0.866 0.255 ;
      LAYER M2 ;
        RECT MASK 1 0.647 0.223 1.09 0.257 ;
        RECT 0.647 0.223 1.09 0.257 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.078 0.647 ;
        RECT MASK 1 -0.042 0.553 1.078 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.078 0.047 ;
        RECT MASK 1 -0.042 -0.047 1.078 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.76 0.454 0.942 0.488 ;
      RECT MASK 1 0.612 0.317 0.646 0.488 ;
      RECT MASK 1 0.612 0.283 0.72 0.317 ;
      RECT MASK 1 0.612 0.132 0.646 0.283 ;
      RECT MASK 1 0.242 0.454 0.572 0.488 ;
      RECT MASK 1 0.538 0.267 0.572 0.454 ;
      RECT MASK 1 0.317 0.243 0.351 0.454 ;
      RECT MASK 1 0.242 0.209 0.351 0.243 ;
      RECT MASK 1 0.242 0.112 0.276 0.209 ;
      RECT MASK 1 0.168 0.317 0.202 0.488 ;
      RECT MASK 1 0.168 0.283 0.276 0.317 ;
      RECT MASK 1 0.168 0.105 0.202 0.283 ;
      RECT MASK 1 0.834 0.186 0.868 0.414 ;
      RECT MASK 1 0.316 0.105 0.424 0.153 ;
      RECT MASK 1 0.76 0.112 0.942 0.146 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.11 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.962 0.55 ;
      RECT 0.074 0.4 0.222 0.45 ;
      RECT 0.37 0.4 0.962 0.45 ;
      RECT 0.814 0.35 0.962 0.4 ;
      RECT 0.222 0.2 0.37 0.25 ;
      RECT 0.074 0.15 0.518 0.2 ;
      RECT 0.666 0.15 0.962 0.2 ;
      RECT 0.074 0.05 0.962 0.15 ;
    LAYER PO ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_ND2B_0P75

MACRO SAEDRVT14_ND2_1P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.666 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.28 0.345 0.31 0.375 ;
        RECT 0.504 0.345 0.534 0.375 ;
      LAYER M2 ;
        RECT MASK 1 0.255 0.343 0.548 0.377 ;
        RECT 0.255 0.343 0.548 0.377 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.102 0.128 0.349 ;
        RECT MASK 1 0.094 0.136 0.128 0.349 ;
        RECT MASK 1 0.398 0.136 0.432 0.349 ;
        RECT MASK 1 0.094 0.102 0.432 0.136 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.201 0.405 0.231 0.435 ;
        RECT 0.585 0.405 0.615 0.435 ;
      LAYER M2 ;
        RECT 0.181 0.403 0.621 0.437 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.708 0.647 ;
        RECT MASK 1 -0.042 0.553 0.708 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.708 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.708 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.086 0.449 0.617 0.483 ;
      RECT MASK 1 0.199 0.21 0.233 0.449 ;
      RECT MASK 1 0.583 0.21 0.617 0.449 ;
      RECT MASK 1 0.199 0.176 0.291 0.21 ;
      RECT MASK 1 0.517 0.176 0.617 0.21 ;
      RECT MASK 1 0.497 0.25 0.543 0.403 ;
      RECT MASK 1 0.273 0.25 0.319 0.403 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.74 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.592 0.55 ;
      RECT 0.074 0.4 0.215 0.45 ;
      RECT 0.303 0.4 0.592 0.45 ;
      RECT 0.074 0.2 0.289 0.25 ;
      RECT 0.377 0.2 0.592 0.25 ;
      RECT 0.074 0.05 0.592 0.2 ;
    LAYER PO ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_ND2_1P5

MACRO SAEDRVT14_NR3_ECO_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.258 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.202 0.276 0.391 ;
        RECT 0.242 0.202 0.276 0.391 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.39 0.202 0.424 0.381 ;
        RECT 0.39 0.202 0.424 0.381 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER VIA1 ;
        RECT 0.594 0.345 0.624 0.375 ;
      LAYER M2 ;
        RECT 0.493 0.343 0.7 0.377 ;
        RECT MASK 1 0.493 0.343 0.7 0.377 ;
    END
  END A3
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.834 0.102 0.868 0.48 ;
        RECT MASK 1 0.834 0.43 0.932 0.48 ;
        RECT MASK 1 0.834 0.152 0.868 0.43 ;
        RECT MASK 1 0.834 0.102 0.932 0.152 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 1.3 0.647 ;
        RECT MASK 1 -0.042 0.553 1.3 0.647 ;
        RECT MASK 1 0.612 0.445 0.646 0.553 ;
        RECT MASK 1 0.76 0.379 0.794 0.553 ;
        RECT MASK 1 1.056 0.451 1.09 0.553 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 1.3 0.047 ;
        RECT MASK 1 0.76 0.047 0.794 0.203 ;
        RECT MASK 1 1.056 0.047 1.09 0.165 ;
        RECT MASK 1 0.094 0.047 0.128 0.16 ;
        RECT MASK 1 0.464 0.047 0.498 0.16 ;
        RECT MASK 1 0.612 0.047 0.646 0.16 ;
        RECT MASK 1 -0.042 -0.047 1.3 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.982 0.088 1.016 0.488 ;
      RECT MASK 1 0.094 0.349 0.128 0.488 ;
      RECT MASK 1 0.094 0.315 0.202 0.349 ;
      RECT MASK 1 0.168 0.154 0.202 0.315 ;
      RECT MASK 1 0.168 0.103 0.389 0.154 ;
      RECT MASK 1 1.13 0.092 1.164 0.484 ;
      RECT MASK 1 0.46 0.445 0.572 0.481 ;
      RECT MASK 1 0.46 0.369 0.498 0.445 ;
      RECT MASK 1 0.168 0.422 0.363 0.472 ;
      RECT MASK 1 0.538 0.363 0.626 0.405 ;
      RECT MASK 1 0.592 0.272 0.626 0.363 ;
      RECT MASK 1 0.908 0.202 0.942 0.374 ;
      RECT MASK 1 0.538 0.087 0.572 0.237 ;
    LAYER M2 ;
      RECT MASK 1 0.133 0.103 1.171 0.137 ;
    LAYER VIA1 ;
      RECT 0.984 0.285 1.014 0.315 ;
      RECT 0.91 0.285 0.94 0.315 ;
      RECT 1.132 0.105 1.162 0.135 ;
      RECT 0.54 0.105 0.57 0.135 ;
      RECT 0.28 0.105 0.31 0.135 ;
    LAYER NWELL ;
      RECT -0.074 0.3 1.332 0.6 ;
    LAYER DIFF ;
      RECT 0.962 0.45 1.11 0.55 ;
      RECT 0.74 0.35 0.888 0.55 ;
      RECT 0.518 0.35 0.666 0.55 ;
      RECT 0.296 0.35 0.444 0.55 ;
      RECT 0.074 0.35 0.222 0.55 ;
      RECT 0.962 0.05 1.11 0.25 ;
      RECT 0.74 0.05 0.888 0.25 ;
      RECT 0.518 0.05 0.666 0.25 ;
      RECT 0.296 0.05 0.444 0.2 ;
      RECT 0.074 0.05 0.222 0.2 ;
    LAYER PO ;
      RECT 1.251 0 1.265 0.6 ;
      RECT 1.177 0 1.191 0.6 ;
      RECT 1.103 0 1.117 0.6 ;
      RECT 1.029 0 1.043 0.6 ;
      RECT 0.955 0 0.969 0.6 ;
      RECT 0.881 0 0.895 0.6 ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_NR3_ECO_1

MACRO SAEDRVT14_AOI21_1P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.74 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.2 0.276 0.348 ;
        RECT 0.242 0.2 0.276 0.348 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.388 0.362 0.422 ;
        RECT MASK 1 0.094 0.158 0.128 0.388 ;
        RECT MASK 1 0.328 0.317 0.362 0.388 ;
        RECT MASK 1 0.328 0.283 0.43 0.317 ;
        RECT 0.094 0.158 0.128 0.422 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.538 0.199 0.572 0.348 ;
        RECT 0.538 0.199 0.572 0.348 ;
    END
  END B
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.458 0.388 0.646 0.422 ;
        RECT MASK 1 0.612 0.15 0.646 0.388 ;
        RECT MASK 1 0.224 0.116 0.646 0.15 ;
        RECT 0.612 0.116 0.646 0.422 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.782 0.647 ;
        RECT MASK 1 -0.042 0.553 0.782 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.782 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.782 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.146 0.462 0.618 0.496 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.814 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.35 0.666 0.55 ;
      RECT 0.155 0.2 0.363 0.25 ;
      RECT 0.074 0.15 0.444 0.2 ;
      RECT 0.074 0.05 0.666 0.15 ;
    LAYER PO ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_AOI21_1P5

MACRO SAEDRVT14_NR2_1P5
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.518 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.242 0.176 0.276 0.338 ;
        RECT MASK 1 0.242 0.176 0.276 0.338 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.094 0.22 0.128 0.488 ;
        RECT MASK 1 0.094 0.454 0.42 0.488 ;
        RECT MASK 1 0.094 0.22 0.128 0.454 ;
        RECT MASK 1 0.386 0.22 0.42 0.454 ;
    END
  END A2
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.234 0.38 0.35 0.414 ;
        RECT MASK 1 0.316 0.15 0.35 0.38 ;
        RECT MASK 1 0.15 0.112 0.388 0.15 ;
        RECT 0.316 0.112 0.35 0.414 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.56 0.647 ;
        RECT MASK 1 -0.042 0.553 0.56 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.56 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.56 0.047 ;
    END
  END VSS
  OBS
    LAYER NWELL ;
      RECT -0.074 0.3 0.592 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.4 0.444 0.55 ;
      RECT 0.074 0.05 0.289 0.25 ;
    LAYER PO ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_NR2_1P5

MACRO SAEDRVT14_NR3_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.814 BY 0.6 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.242 0.199 0.276 0.445 ;
        RECT 0.242 0.199 0.276 0.445 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.168 0.199 0.202 0.505 ;
        RECT MASK 1 0.168 0.199 0.202 0.505 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.094 0.197 0.128 0.458 ;
        RECT 0.094 0.197 0.128 0.458 ;
    END
  END A3
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT MASK 1 0.612 0.099 0.646 0.507 ;
        RECT 0.612 0.099 0.646 0.507 ;
    END
  END X
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M1 ;
        RECT -0.042 0.553 0.856 0.647 ;
        RECT MASK 1 -0.042 0.553 0.856 0.647 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -0.042 -0.047 0.856 0.047 ;
        RECT MASK 1 -0.042 -0.047 0.856 0.047 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT MASK 1 0.442 0.454 0.572 0.488 ;
      RECT MASK 1 0.538 0.146 0.572 0.454 ;
      RECT MASK 1 0.442 0.112 0.572 0.146 ;
      RECT MASK 1 0.316 0.316 0.35 0.488 ;
      RECT MASK 1 0.427 0.316 0.461 0.414 ;
      RECT MASK 1 0.316 0.282 0.461 0.316 ;
      RECT MASK 1 0.427 0.186 0.461 0.282 ;
      RECT MASK 1 0.316 0.146 0.35 0.282 ;
      RECT MASK 1 0.146 0.112 0.35 0.146 ;
    LAYER NWELL ;
      RECT -0.074 0.3 0.888 0.6 ;
    LAYER DIFF ;
      RECT 0.074 0.45 0.74 0.55 ;
      RECT 0.074 0.35 0.37 0.45 ;
      RECT 0.518 0.35 0.74 0.45 ;
      RECT 0.074 0.2 0.289 0.25 ;
      RECT 0.37 0.2 0.74 0.25 ;
      RECT 0.074 0.05 0.74 0.2 ;
    LAYER PO ;
      RECT 0.807 0 0.821 0.6 ;
      RECT 0.733 0 0.747 0.6 ;
      RECT 0.659 0 0.673 0.6 ;
      RECT 0.585 0 0.599 0.6 ;
      RECT 0.511 0 0.525 0.6 ;
      RECT 0.437 0 0.451 0.6 ;
      RECT 0.363 0 0.377 0.6 ;
      RECT 0.289 0 0.303 0.6 ;
      RECT 0.215 0 0.229 0.6 ;
      RECT 0.141 0 0.155 0.6 ;
      RECT 0.067 0 0.081 0.6 ;
      RECT -0.007 0 0.007 0.6 ;
  END
END SAEDRVT14_NR3_2

END LIBRARY
