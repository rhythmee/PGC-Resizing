VERSION 5.8 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.001 ;

PROPERTYDEFINITIONS
  MACRO expanded_util REAL ;
  MACRO previous_effective_target_usage REAL ;
END PROPERTYDEFINITIONS

LAYER NWELL
  TYPE MASTERSLICE ;
END NWELL

LAYER PO
  TYPE MASTERSLICE ;
END PO

LAYER CO
  TYPE CUT ;
END CO

LAYER M1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.152 ;
  WIDTH 0.05 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.05 WRONGDIRECTION ;" ;
END M1

LAYER VIA1
  TYPE CUT ;
END VIA1

LAYER M2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.152 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M2

LAYER VIA2
  TYPE CUT ;
END VIA2

LAYER M3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.304 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M3

LAYER VIA3
  TYPE CUT ;
END VIA3

LAYER M4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.304 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M4

LAYER VIA4
  TYPE CUT ;
END VIA4

LAYER M5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.608 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M5

LAYER VIA5
  TYPE CUT ;
END VIA5

LAYER M6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.608 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M6

LAYER VIA6
  TYPE CUT ;
END VIA6

LAYER M7
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 1.216 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M7

LAYER VIA7
  TYPE CUT ;
END VIA7

LAYER M8
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 1.216 ;
  WIDTH 0.056 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.056 WRONGDIRECTION ;" ;
END M8

LAYER VIA8
  TYPE CUT ;
END VIA8

LAYER M9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 2.432 ;
  WIDTH 0.16 ;
  PROPERTY LEF58_WIDTH "WIDTH 0.16 WRONGDIRECTION ;" ;
END M9

LAYER VIARDL
  TYPE CUT ;
END VIARDL

LAYER MRDL
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 4.864 ;
  WIDTH 2 ;
  PROPERTY LEF58_WIDTH "WIDTH 2 WRONGDIRECTION ;" ;
END MRDL

LAYER DNW
  TYPE MASTERSLICE ;
END DNW

LAYER DIFF
  TYPE MASTERSLICE ;
END DIFF

LAYER PIMP
  TYPE MASTERSLICE ;
END PIMP

LAYER NIMP
  TYPE MASTERSLICE ;
END NIMP

LAYER DIFF_18
  TYPE MASTERSLICE ;
END DIFF_18

LAYER PAD
  TYPE MASTERSLICE ;
END PAD

LAYER ESD_25
  TYPE MASTERSLICE ;
END ESD_25

LAYER SBLK
  TYPE MASTERSLICE ;
END SBLK

LAYER HVTIMP
  TYPE MASTERSLICE ;
END HVTIMP

LAYER LVTIMP
  TYPE MASTERSLICE ;
END LVTIMP

LAYER M1PIN
  TYPE MASTERSLICE ;
END M1PIN

LAYER M2PIN
  TYPE MASTERSLICE ;
END M2PIN

LAYER M3PIN
  TYPE MASTERSLICE ;
END M3PIN

LAYER M4PIN
  TYPE MASTERSLICE ;
END M4PIN

LAYER M5PIN
  TYPE MASTERSLICE ;
END M5PIN

LAYER M6PIN
  TYPE MASTERSLICE ;
END M6PIN

LAYER M7PIN
  TYPE MASTERSLICE ;
END M7PIN

LAYER M8PIN
  TYPE MASTERSLICE ;
END M8PIN

LAYER M9PIN
  TYPE MASTERSLICE ;
END M9PIN

LAYER MRDL9PIN
  TYPE MASTERSLICE ;
END MRDL9PIN

LAYER HOTNWL
  TYPE MASTERSLICE ;
END HOTNWL

LAYER DIOD
  TYPE MASTERSLICE ;
END DIOD

LAYER BJTDMY
  TYPE MASTERSLICE ;
END BJTDMY

LAYER RNW
  TYPE MASTERSLICE ;
END RNW

LAYER RMARK
  TYPE MASTERSLICE ;
END RMARK

LAYER prBoundary
  TYPE MASTERSLICE ;
END prBoundary

LAYER LOGO
  TYPE MASTERSLICE ;
END LOGO

LAYER IP
  TYPE MASTERSLICE ;
END IP

LAYER RM1
  TYPE MASTERSLICE ;
END RM1

LAYER RM2
  TYPE MASTERSLICE ;
END RM2

LAYER RM3
  TYPE MASTERSLICE ;
END RM3

LAYER RM4
  TYPE MASTERSLICE ;
END RM4

LAYER RM5
  TYPE MASTERSLICE ;
END RM5

LAYER RM6
  TYPE MASTERSLICE ;
END RM6

LAYER RM7
  TYPE MASTERSLICE ;
END RM7

LAYER RM8
  TYPE MASTERSLICE ;
END RM8

LAYER RM9
  TYPE MASTERSLICE ;
END RM9

LAYER DM1EXCL
  TYPE MASTERSLICE ;
END DM1EXCL

LAYER DM2EXCL
  TYPE MASTERSLICE ;
END DM2EXCL

LAYER DM3EXCL
  TYPE MASTERSLICE ;
END DM3EXCL

LAYER DM4EXCL
  TYPE MASTERSLICE ;
END DM4EXCL

LAYER DM5EXCL
  TYPE MASTERSLICE ;
END DM5EXCL

LAYER DM6EXCL
  TYPE MASTERSLICE ;
END DM6EXCL

LAYER DM7EXCL
  TYPE MASTERSLICE ;
END DM7EXCL

LAYER DM8EXCL
  TYPE MASTERSLICE ;
END DM8EXCL

LAYER DM9EXCL
  TYPE MASTERSLICE ;
END DM9EXCL

LAYER DIFF_25
  TYPE MASTERSLICE ;
END DIFF_25

LAYER DIFF_FM
  TYPE MASTERSLICE ;
END DIFF_FM

LAYER PO_FM
  TYPE MASTERSLICE ;
END PO_FM

VIA VIA12SQ_C
  LAYER M1 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA12SQ_C

VIA VIA12BAR_C
  LAYER M1 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M2 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA12BAR_C

VIA VIA12LG_C
  LAYER M1 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA12LG_C

VIA VIA12SQ
  LAYER M1 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA1 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA12SQ

VIA VIA12BAR
  LAYER M1 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA1 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA12BAR

VIA VIA12LG
  LAYER M1 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA12LG

VIA VIA23SQ_C
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA23SQ_C

VIA VIA23BAR_C
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M3 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA23BAR_C

VIA VIA23LG_C
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA23LG_C

VIA VIA23SQ
  LAYER M2 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA2 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA23SQ

VIA VIA23BAR
  LAYER M2 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA2 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA23BAR

VIA VIA23LG
  LAYER M2 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA23LG

VIA VIA34SQ_C
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA34SQ_C

VIA VIA34BAR_C
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M4 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA34BAR_C

VIA VIA34LG_C
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA34LG_C

VIA VIA34SQ
  LAYER M3 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA3 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA34SQ

VIA VIA34BAR
  LAYER M3 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA3 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA34BAR

VIA VIA34LG
  LAYER M3 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA34LG

VIA VIA45SQ_C
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA45SQ_C

VIA VIA45BAR_C
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA4 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M5 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA45BAR_C

VIA VIA45LG_C
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA45LG_C

VIA VIA45SQ
  LAYER M4 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA4 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M5 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA45SQ

VIA VIA45BAR
  LAYER M4 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA4 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA45BAR

VIA VIA45LG
  LAYER M4 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA45LG

VIA VIA56SQ_C
  LAYER M5 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA56SQ_C

VIA VIA56BAR_C
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M6 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA56BAR_C

VIA VIA56LG_C
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA56LG_C

VIA VIA56SQ
  LAYER M5 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA5 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA56SQ

VIA VIA56BAR
  LAYER M5 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA5 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA56BAR

VIA VIA56LG
  LAYER M5 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA56LG

VIA VIA67SQ_C
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA6 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M7 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA67SQ_C

VIA VIA67BAR_C
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA6 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M7 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA67BAR_C

VIA VIA67LG_C
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA67LG_C

VIA VIA67SQ
  LAYER M6 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA6 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M7 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA67SQ

VIA VIA67BAR
  LAYER M6 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA6 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA67BAR

VIA VIA67LG
  LAYER M6 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA67LG

VIA VIA78SQ_C
  LAYER M7 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA7 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M8 ;
    RECT -0.03 -0.055 0.03 0.055 ;
END VIA78SQ_C

VIA VIA78BAR_C
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA7 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M8 ;
    RECT -0.03 -0.08 0.03 0.08 ;
END VIA78BAR_C

VIA VIA78LG_C
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA7 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M8 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA78LG_C

VIA VIA78SQ
  LAYER M7 ;
    RECT -0.055 -0.03 0.055 0.03 ;
  LAYER VIA7 ;
    RECT -0.025 -0.025 0.025 0.025 ;
  LAYER M8 ;
    RECT -0.055 -0.03 0.055 0.03 ;
END VIA78SQ

VIA VIA78BAR
  LAYER M7 ;
    RECT -0.055 -0.055 0.055 0.055 ;
  LAYER VIA7 ;
    RECT -0.025 -0.05 0.025 0.05 ;
  LAYER M8 ;
    RECT -0.055 -0.055 0.055 0.055 ;
END VIA78BAR

VIA VIA78LG
  LAYER M7 ;
    RECT -0.08 -0.055 0.08 0.055 ;
  LAYER VIA7 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M8 ;
    RECT -0.08 -0.055 0.08 0.055 ;
END VIA78LG

VIA VIA89_C
  LAYER M8 ;
    RECT -0.095 -0.08 0.095 0.08 ;
  LAYER VIA8 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M9 ;
    RECT -0.08 -0.095 0.08 0.095 ;
END VIA89_C

VIA VIA89
  LAYER M8 ;
    RECT -0.095 -0.08 0.095 0.08 ;
  LAYER VIA8 ;
    RECT -0.065 -0.065 0.065 0.065 ;
  LAYER M9 ;
    RECT -0.095 -0.08 0.095 0.08 ;
END VIA89

VIA VIA9RDL
  LAYER M9 ;
    RECT -1.5 -1.5 1.5 1.5 ;
  LAYER VIARDL ;
    RECT -1 -1 1 1 ;
  LAYER MRDL ;
    RECT -1.5 -1.5 1.5 1.5 ;
END VIA9RDL

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.152 BY 1.672 ;
END unit

MACRO DFFX1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.952 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.684 0.401 0.726 ;
      LAYER M1 ;
        RECT 0.249 0.68 0.421 0.73 ;
        RECT 0.249 0.553 0.359 0.68 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 ;
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 1.53 0.705 1.572 ;
      LAYER M1 ;
        RECT 0.553 1.424 0.725 1.576 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.323 0.195 3.365 0.237 ;
        RECT 3.323 0.287 3.365 0.329 ;
        RECT 3.323 0.932 3.365 0.974 ;
        RECT 3.323 1.024 3.365 1.066 ;
        RECT 3.323 1.116 3.365 1.158 ;
        RECT 3.323 1.208 3.365 1.25 ;
        RECT 3.323 1.3 3.365 1.342 ;
        RECT 3.323 1.392 3.365 1.434 ;
        RECT 3.323 1.484 3.365 1.526 ;
      LAYER M1 ;
        RECT 3.593 1.009 3.703 1.119 ;
        RECT 3.319 0.854 3.369 1.546 ;
        RECT 3.653 0.854 3.703 1.009 ;
        RECT 3.319 0.804 3.703 0.854 ;
        RECT 3.653 0.359 3.703 0.804 ;
        RECT 3.319 0.309 3.703 0.359 ;
        RECT 3.319 0.148 3.369 0.309 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.627 0.158 3.669 0.2 ;
        RECT 3.627 1.3 3.669 1.342 ;
        RECT 3.627 1.392 3.669 1.434 ;
        RECT 3.627 1.484 3.669 1.526 ;
      LAYER M1 ;
        RECT 3.623 1.271 3.673 1.546 ;
        RECT 3.623 1.221 3.856 1.271 ;
        RECT 3.745 1.161 3.856 1.221 ;
        RECT 3.805 0.204 3.855 1.161 ;
        RECT 3.607 0.154 3.855 0.204 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.062 0.325 1.104 ;
        RECT 3.475 1.072 3.517 1.114 ;
        RECT 0.739 1.108 0.781 1.15 ;
        RECT 0.891 1.122 0.933 1.164 ;
        RECT 0.283 1.154 0.325 1.196 ;
        RECT 3.475 1.164 3.517 1.206 ;
        RECT 0.739 1.2 0.781 1.242 ;
        RECT 0.891 1.214 0.933 1.256 ;
        RECT 3.475 1.256 3.517 1.298 ;
        RECT 1.803 1.282 1.845 1.324 ;
        RECT 1.955 1.282 1.997 1.324 ;
        RECT 0.739 1.292 0.781 1.334 ;
        RECT 0.891 1.306 0.933 1.348 ;
        RECT 2.715 1.312 2.757 1.354 ;
        RECT 3.171 1.312 3.213 1.354 ;
        RECT 3.475 1.348 3.517 1.39 ;
        RECT 0.891 1.398 0.933 1.44 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
        RECT 3.095 1.651 3.137 1.693 ;
        RECT 3.247 1.651 3.289 1.693 ;
        RECT 3.399 1.651 3.441 1.693 ;
        RECT 3.551 1.651 3.593 1.693 ;
        RECT 3.703 1.651 3.745 1.693 ;
        RECT 3.855 1.651 3.897 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 3.952 1.702 ;
        RECT 2.639 1.358 2.689 1.642 ;
        RECT 3.207 1.358 3.257 1.642 ;
        RECT 0.887 1.354 0.937 1.642 ;
        RECT 1.975 1.328 2.025 1.642 ;
        RECT 2.639 1.308 2.777 1.358 ;
        RECT 3.149 1.308 3.257 1.358 ;
        RECT 0.279 1.033 0.329 1.642 ;
        RECT 3.471 0.947 3.521 1.642 ;
        RECT 0.735 1.304 0.937 1.354 ;
        RECT 1.782 1.278 2.025 1.328 ;
        RECT 0.735 1.088 0.785 1.304 ;
        RECT 0.887 1.101 0.937 1.304 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 3.399 -0.021 3.441 0.021 ;
        RECT 3.551 -0.021 3.593 0.021 ;
        RECT 3.703 -0.021 3.745 0.021 ;
        RECT 3.855 -0.021 3.897 0.021 ;
        RECT 3.475 0.158 3.517 0.2 ;
        RECT 0.739 0.2 0.781 0.242 ;
        RECT 1.955 0.203 1.997 0.245 ;
        RECT 1.803 0.219 1.845 0.261 ;
        RECT 0.891 0.275 0.933 0.317 ;
        RECT 1.803 0.311 1.845 0.353 ;
        RECT 2.715 0.334 2.757 0.376 ;
        RECT 3.171 0.334 3.213 0.376 ;
        RECT 0.283 0.344 0.325 0.386 ;
        RECT 0.739 0.388 0.781 0.43 ;
        RECT 0.891 0.388 0.933 0.43 ;
      LAYER M1 ;
        RECT 2.695 0.33 3.233 0.38 ;
        RECT 1.799 0.249 1.849 0.373 ;
        RECT 0.735 0.246 0.785 0.45 ;
        RECT 0.887 0.246 0.937 0.45 ;
        RECT 1.799 0.199 2.024 0.249 ;
        RECT 0.586 0.196 0.937 0.246 ;
        RECT 0.279 0.03 0.329 0.419 ;
        RECT 3.167 0.03 3.217 0.33 ;
        RECT 3.471 0.03 3.521 0.22 ;
        RECT 1.799 0.03 1.849 0.199 ;
        RECT 0.586 0.03 0.636 0.196 ;
        RECT 0 -0.03 3.952 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 1.195 0.319 1.237 0.361 ;
      RECT 1.347 0.375 1.389 0.417 ;
      RECT 1.727 0.762 1.769 0.804 ;
      RECT 1.879 1.522 1.921 1.564 ;
      RECT 1.195 1.252 1.237 1.294 ;
      RECT 1.043 0.506 1.085 0.548 ;
      RECT 0.435 1.062 0.477 1.104 ;
      RECT 1.043 0.414 1.085 0.456 ;
      RECT 0.435 1.154 0.477 1.196 ;
      RECT 0.435 1.062 0.477 1.104 ;
      RECT 2.107 1.199 2.149 1.241 ;
      RECT 2.107 1.291 2.149 1.333 ;
      RECT 2.867 1.212 2.909 1.254 ;
      RECT 1.499 1.162 1.541 1.204 ;
      RECT 1.347 1.16 1.389 1.202 ;
      RECT 1.119 1.53 1.161 1.572 ;
      RECT 1.727 1.482 1.769 1.524 ;
      RECT 0.587 0.76 0.629 0.802 ;
      RECT 2.031 0.644 2.073 0.686 ;
      RECT 2.259 1.107 2.301 1.149 ;
      RECT 3.095 1.525 3.137 1.567 ;
      RECT 2.183 1.526 2.225 1.568 ;
      RECT 1.271 1.49 1.313 1.532 ;
      RECT 2.791 1.525 2.833 1.567 ;
      RECT 3.551 0.608 3.593 0.65 ;
      RECT 2.639 0.703 2.681 0.745 ;
      RECT 2.867 0.442 2.909 0.484 ;
      RECT 2.411 0.49 2.453 0.532 ;
      RECT 2.183 0.644 2.225 0.686 ;
      RECT 2.791 0.12 2.833 0.162 ;
      RECT 2.335 0.18 2.377 0.222 ;
      RECT 1.727 0.544 1.769 0.586 ;
      RECT 1.499 0.438 1.541 0.48 ;
      RECT 1.423 0.1 1.465 0.142 ;
      RECT 2.943 0.608 2.985 0.65 ;
      RECT 1.575 1.005 1.617 1.047 ;
      RECT 0.815 0.1 0.857 0.142 ;
      RECT 1.119 0.649 1.161 0.691 ;
      RECT 0.435 0.492 0.477 0.534 ;
      RECT 1.195 1.16 1.237 1.202 ;
      RECT 2.335 1.526 2.377 1.568 ;
      RECT 1.043 0.852 1.085 0.894 ;
      RECT 2.259 0.391 2.301 0.433 ;
      RECT 3.399 0.608 3.441 0.65 ;
      RECT 2.563 0.982 2.605 1.024 ;
      RECT 1.043 0.76 1.085 0.802 ;
      RECT 0.815 0.622 0.857 0.664 ;
      RECT 2.259 1.291 2.301 1.333 ;
      RECT 0.435 1.154 0.477 1.196 ;
      RECT 2.411 1.103 2.453 1.145 ;
      RECT 2.107 0.424 2.149 0.466 ;
      RECT 0.967 0.622 1.009 0.664 ;
      RECT 1.347 1.252 1.389 1.294 ;
      RECT 2.563 0.542 2.605 0.584 ;
      RECT 1.879 0.544 1.921 0.586 ;
      RECT 1.423 1.503 1.465 1.545 ;
      RECT 2.259 1.199 2.301 1.241 ;
      RECT 0.587 0.442 0.629 0.484 ;
      RECT 0.587 0.442 0.629 0.484 ;
      RECT 1.271 0.1 1.313 0.142 ;
      RECT 0.587 0.442 0.629 0.484 ;
      RECT 1.347 0.375 1.389 0.417 ;
      RECT 1.347 0.375 1.389 0.417 ;
      RECT 1.195 0.319 1.237 0.361 ;
      RECT 1.195 0.319 1.237 0.361 ;
      RECT 0.587 0.852 0.629 0.894 ;
      RECT 3.095 0.713 3.137 0.755 ;
    LAYER M1 ;
      RECT 1.191 0.299 1.281 0.381 ;
      RECT 0.431 0.988 1.265 1.038 ;
      RECT 1.191 1.038 1.241 1.314 ;
      RECT 1.215 0.381 1.265 0.988 ;
      RECT 0.431 0.779 0.521 0.829 ;
      RECT 0.431 0.579 0.521 0.629 ;
      RECT 0.431 1.038 0.481 1.216 ;
      RECT 0.431 0.829 0.481 0.988 ;
      RECT 0.431 0.455 0.481 0.579 ;
      RECT 0.471 0.629 0.521 0.779 ;
      RECT 2.115 0.23 2.837 0.28 ;
      RECT 2.787 0.088 2.837 0.23 ;
      RECT 1.964 0.314 2.165 0.364 ;
      RECT 1.707 0.54 2.014 0.59 ;
      RECT 2.315 0.178 2.397 0.23 ;
      RECT 2.115 0.28 2.165 0.314 ;
      RECT 1.964 0.364 2.014 0.54 ;
      RECT 1.343 0.64 2.093 0.69 ;
      RECT 1.343 0.434 1.561 0.484 ;
      RECT 1.343 1.158 1.561 1.208 ;
      RECT 1.343 0.355 1.393 0.434 ;
      RECT 1.343 1.208 1.393 1.314 ;
      RECT 1.343 0.69 1.393 1.158 ;
      RECT 1.343 0.484 1.393 0.64 ;
      RECT 3.207 0.704 3.597 0.754 ;
      RECT 2.407 0.438 3.597 0.488 ;
      RECT 3.547 0.488 3.597 0.704 ;
      RECT 2.619 0.699 2.76 0.749 ;
      RECT 2.847 1.208 3.257 1.258 ;
      RECT 2.407 0.488 2.457 1.165 ;
      RECT 2.71 0.488 2.76 0.699 ;
      RECT 3.207 0.754 3.257 1.208 ;
      RECT 1.707 0.758 2.229 0.808 ;
      RECT 2.179 0.587 2.229 0.758 ;
      RECT 1.55 1.001 2.345 1.051 ;
      RECT 2.255 0.371 2.305 0.42 ;
      RECT 2.072 0.42 2.345 0.47 ;
      RECT 2.103 1.166 2.153 1.308 ;
      RECT 2.103 1.308 2.305 1.358 ;
      RECT 2.295 0.47 2.345 1.001 ;
      RECT 2.255 1.051 2.305 1.308 ;
      RECT 2.824 0.604 3.461 0.654 ;
      RECT 2.519 0.538 2.649 0.588 ;
      RECT 2.824 1.028 2.874 1.029 ;
      RECT 2.824 0.654 2.874 0.978 ;
      RECT 2.542 1.027 2.874 1.028 ;
      RECT 2.519 0.588 2.569 0.978 ;
      RECT 2.519 0.978 2.874 1.027 ;
      RECT 2.77 1.521 3.157 1.571 ;
      RECT 1.419 1.478 1.789 1.528 ;
      RECT 1.419 1.528 1.469 1.565 ;
      RECT 1.099 1.526 1.317 1.576 ;
      RECT 1.875 1.428 1.925 1.584 ;
      RECT 1.267 1.428 1.317 1.526 ;
      RECT 1.267 1.378 1.925 1.428 ;
      RECT 0.583 0.618 1.029 0.668 ;
      RECT 0.583 0.668 0.633 0.914 ;
      RECT 0.583 0.422 0.633 0.618 ;
      RECT 1.039 0.518 1.165 0.568 ;
      RECT 1.039 0.768 1.089 0.914 ;
      RECT 1.039 0.718 1.165 0.768 ;
      RECT 1.039 0.394 1.089 0.518 ;
      RECT 1.115 0.568 1.165 0.718 ;
      RECT 2.934 0.709 3.157 0.759 ;
      RECT 2.355 1.272 2.581 1.322 ;
      RECT 2.163 1.522 2.405 1.572 ;
      RECT 2.355 1.322 2.405 1.522 ;
      RECT 2.531 1.149 2.581 1.272 ;
      RECT 2.934 0.759 2.984 1.099 ;
      RECT 2.531 1.099 2.984 1.149 ;
      RECT 0.795 0.096 1.491 0.146 ;
    LAYER PO ;
      RECT 3.101 1.012 3.131 1.606 ;
      RECT 2.341 0.068 2.371 0.622 ;
      RECT 0.061 0.066 0.091 1.606 ;
      RECT 0.365 0.068 0.395 1.606 ;
      RECT 0.213 0.066 0.243 1.606 ;
      RECT 1.733 0.73 1.763 1.606 ;
      RECT 1.125 0.068 1.155 1.606 ;
      RECT 3.253 0.068 3.283 1.606 ;
      RECT 3.709 0.068 3.739 1.606 ;
      RECT 2.949 0.068 2.979 1.606 ;
      RECT 1.885 0.068 1.915 1.606 ;
      RECT 0.669 0.068 0.699 1.606 ;
      RECT 2.037 0.068 2.067 1.606 ;
      RECT 1.581 0.068 1.611 1.606 ;
      RECT 0.821 0.068 0.851 1.606 ;
      RECT 2.493 0.068 2.523 1.606 ;
      RECT 2.189 0.068 2.219 1.606 ;
      RECT 2.797 0.068 2.827 1.606 ;
      RECT 3.557 0.068 3.587 1.606 ;
      RECT 1.429 0.068 1.459 1.606 ;
      RECT 2.645 0.068 2.675 1.606 ;
      RECT 0.973 0.068 1.003 1.606 ;
      RECT 3.405 0.068 3.435 1.606 ;
      RECT 0.517 0.068 0.547 1.606 ;
      RECT 1.277 0.068 1.307 0.542 ;
      RECT 3.861 0.068 3.891 1.606 ;
      RECT 1.277 0.99 1.307 1.606 ;
      RECT 3.101 0.068 3.131 0.787 ;
      RECT 1.733 0.068 1.763 0.618 ;
      RECT 2.341 0.882 2.371 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 4.067 1.773 ;
  END
END DFFX1_RVT

MACRO DFFARX1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 4.256 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.684 0.401 0.726 ;
      LAYER M1 ;
        RECT 0.249 0.68 0.421 0.73 ;
        RECT 0.249 0.553 0.359 0.68 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 ;
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 1.53 0.705 1.572 ;
      LAYER M1 ;
        RECT 0.553 1.424 0.725 1.576 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 2.791 0.124 2.833 0.166 ;
        RECT 1.727 0.138 1.769 0.18 ;
      LAYER M1 ;
        RECT 1.723 0.144 1.879 0.223 ;
        RECT 2.771 0.144 2.853 0.18 ;
        RECT 1.723 0.094 2.853 0.144 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0441 ;
  END RSTB
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.627 0.195 3.669 0.237 ;
        RECT 3.627 0.287 3.669 0.329 ;
        RECT 3.627 0.932 3.669 0.974 ;
        RECT 3.627 1.024 3.669 1.066 ;
        RECT 3.627 1.116 3.669 1.158 ;
        RECT 3.627 1.208 3.669 1.25 ;
        RECT 3.627 1.3 3.669 1.342 ;
        RECT 3.627 1.392 3.669 1.434 ;
        RECT 3.627 1.484 3.669 1.526 ;
      LAYER M1 ;
        RECT 3.897 1.009 4.007 1.119 ;
        RECT 3.623 0.854 3.673 1.546 ;
        RECT 3.957 0.854 4.007 1.009 ;
        RECT 3.623 0.804 4.007 0.854 ;
        RECT 3.957 0.359 4.007 0.804 ;
        RECT 3.623 0.309 4.007 0.359 ;
        RECT 3.623 0.148 3.673 0.309 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.931 0.158 3.973 0.2 ;
        RECT 3.931 1.3 3.973 1.342 ;
        RECT 3.931 1.392 3.973 1.434 ;
        RECT 3.931 1.484 3.973 1.526 ;
      LAYER M1 ;
        RECT 3.927 1.271 3.977 1.546 ;
        RECT 3.927 1.221 4.16 1.271 ;
        RECT 4.05 1.161 4.16 1.221 ;
        RECT 4.109 0.204 4.159 1.161 ;
        RECT 3.911 0.154 4.159 0.204 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.062 0.325 1.104 ;
        RECT 3.779 1.072 3.821 1.114 ;
        RECT 0.739 1.118 0.781 1.16 ;
        RECT 0.891 1.132 0.933 1.174 ;
        RECT 0.283 1.154 0.325 1.196 ;
        RECT 3.779 1.164 3.821 1.206 ;
        RECT 0.739 1.21 0.781 1.252 ;
        RECT 0.891 1.224 0.933 1.266 ;
        RECT 3.779 1.256 3.821 1.298 ;
        RECT 1.955 1.282 1.997 1.324 ;
        RECT 2.107 1.282 2.149 1.324 ;
        RECT 0.739 1.302 0.781 1.344 ;
        RECT 2.867 1.312 2.909 1.354 ;
        RECT 3.475 1.312 3.517 1.354 ;
        RECT 0.891 1.316 0.933 1.358 ;
        RECT 3.779 1.348 3.821 1.39 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
        RECT 3.095 1.651 3.137 1.693 ;
        RECT 3.247 1.651 3.289 1.693 ;
        RECT 3.399 1.651 3.441 1.693 ;
        RECT 3.551 1.651 3.593 1.693 ;
        RECT 3.703 1.651 3.745 1.693 ;
        RECT 3.855 1.651 3.897 1.693 ;
        RECT 4.007 1.651 4.049 1.693 ;
        RECT 4.159 1.651 4.201 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 4.256 1.702 ;
        RECT 0.887 1.364 0.937 1.642 ;
        RECT 3.511 1.358 3.561 1.642 ;
        RECT 2.127 1.328 2.177 1.642 ;
        RECT 0.279 1.033 0.329 1.642 ;
        RECT 3.775 0.947 3.825 1.642 ;
        RECT 0.735 1.314 0.937 1.364 ;
        RECT 2.834 1.308 3.561 1.358 ;
        RECT 1.934 1.278 2.177 1.328 ;
        RECT 0.735 1.098 0.785 1.314 ;
        RECT 0.887 1.111 0.937 1.314 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 3.399 -0.021 3.441 0.021 ;
        RECT 3.551 -0.021 3.593 0.021 ;
        RECT 3.703 -0.021 3.745 0.021 ;
        RECT 3.855 -0.021 3.897 0.021 ;
        RECT 4.007 -0.021 4.049 0.021 ;
        RECT 4.159 -0.021 4.201 0.021 ;
        RECT 3.779 0.158 3.821 0.2 ;
        RECT 0.739 0.2 0.781 0.242 ;
        RECT 2.107 0.203 2.149 0.245 ;
        RECT 0.891 0.275 0.933 0.317 ;
        RECT 1.955 0.307 1.997 0.349 ;
        RECT 3.019 0.334 3.061 0.376 ;
        RECT 3.475 0.334 3.517 0.376 ;
        RECT 0.283 0.344 0.325 0.386 ;
        RECT 0.739 0.388 0.781 0.43 ;
        RECT 0.891 0.388 0.933 0.43 ;
        RECT 1.955 0.399 1.997 0.441 ;
      LAYER M1 ;
        RECT 1.951 0.337 2.001 0.461 ;
        RECT 2.999 0.33 3.537 0.38 ;
        RECT 1.541 0.287 2.001 0.337 ;
        RECT 1.951 0.249 2.001 0.287 ;
        RECT 0.735 0.246 0.785 0.45 ;
        RECT 0.887 0.246 0.937 0.45 ;
        RECT 1.951 0.199 2.176 0.249 ;
        RECT 0.586 0.196 0.937 0.246 ;
        RECT 0.279 0.03 0.329 0.419 ;
        RECT 3.471 0.03 3.521 0.33 ;
        RECT 1.541 0.03 1.591 0.287 ;
        RECT 3.775 0.03 3.825 0.22 ;
        RECT 0.586 0.03 0.636 0.196 ;
        RECT 0 -0.03 4.256 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 2.715 0.982 2.757 1.024 ;
      RECT 1.043 0.76 1.085 0.802 ;
      RECT 0.815 0.622 0.857 0.664 ;
      RECT 2.411 1.291 2.453 1.333 ;
      RECT 0.435 1.154 0.477 1.196 ;
      RECT 2.563 1.103 2.605 1.145 ;
      RECT 3.171 1.212 3.213 1.254 ;
      RECT 0.967 0.622 1.009 0.664 ;
      RECT 1.195 0.319 1.237 0.361 ;
      RECT 1.347 0.375 1.389 0.417 ;
      RECT 1.879 0.79 1.921 0.832 ;
      RECT 3.171 0.442 3.213 0.484 ;
      RECT 0.587 0.442 0.629 0.484 ;
      RECT 0.587 0.442 0.629 0.484 ;
      RECT 0.587 0.442 0.629 0.484 ;
      RECT 1.347 0.375 1.389 0.417 ;
      RECT 1.347 0.375 1.389 0.417 ;
      RECT 1.195 0.319 1.237 0.361 ;
      RECT 1.195 0.319 1.237 0.361 ;
      RECT 0.587 0.852 0.629 0.894 ;
      RECT 0.435 1.154 0.477 1.196 ;
      RECT 0.435 1.062 0.477 1.104 ;
      RECT 3.019 0.982 3.061 1.024 ;
      RECT 2.031 1.492 2.073 1.534 ;
      RECT 1.195 1.252 1.237 1.294 ;
      RECT 1.043 0.506 1.085 0.548 ;
      RECT 0.435 1.062 0.477 1.104 ;
      RECT 1.043 0.414 1.085 0.456 ;
      RECT 3.399 0.713 3.441 0.755 ;
      RECT 3.247 0.608 3.289 0.65 ;
      RECT 1.651 1.162 1.693 1.204 ;
      RECT 1.347 1.16 1.389 1.202 ;
      RECT 0.815 0.1 0.857 0.142 ;
      RECT 1.879 1.482 1.921 1.524 ;
      RECT 0.587 0.76 0.629 0.802 ;
      RECT 2.183 0.672 2.225 0.714 ;
      RECT 2.411 1.107 2.453 1.149 ;
      RECT 2.259 1.282 2.301 1.324 ;
      RECT 2.335 1.532 2.377 1.574 ;
      RECT 1.271 1.49 1.313 1.532 ;
      RECT 3.095 1.433 3.137 1.475 ;
      RECT 1.499 1.282 1.541 1.324 ;
      RECT 3.855 0.608 3.897 0.65 ;
      RECT 2.943 0.77 2.985 0.812 ;
      RECT 2.563 0.49 2.605 0.532 ;
      RECT 3.095 0.172 3.137 0.214 ;
      RECT 2.487 0.218 2.529 0.26 ;
      RECT 1.879 0.572 1.921 0.614 ;
      RECT 1.499 0.438 1.541 0.48 ;
      RECT 2.335 0.641 2.377 0.683 ;
      RECT 1.575 1.005 1.617 1.047 ;
      RECT 1.803 1.282 1.845 1.324 ;
      RECT 1.119 0.649 1.161 0.691 ;
      RECT 0.435 0.492 0.477 0.534 ;
      RECT 1.271 0.1 1.313 0.142 ;
      RECT 1.119 1.53 1.161 1.572 ;
      RECT 1.423 0.1 1.465 0.142 ;
      RECT 2.259 1.164 2.301 1.206 ;
      RECT 1.043 0.852 1.085 0.894 ;
      RECT 2.411 0.391 2.453 0.433 ;
      RECT 3.703 0.608 3.745 0.65 ;
      RECT 3.399 1.432 3.441 1.474 ;
      RECT 1.195 1.16 1.237 1.202 ;
      RECT 2.487 1.532 2.529 1.574 ;
      RECT 2.259 0.424 2.301 0.466 ;
      RECT 1.347 1.252 1.389 1.294 ;
      RECT 2.715 0.542 2.757 0.584 ;
      RECT 2.031 0.572 2.073 0.614 ;
      RECT 1.423 1.503 1.465 1.545 ;
      RECT 2.411 1.199 2.453 1.241 ;
    LAYER M1 ;
      RECT 1.191 0.299 1.281 0.381 ;
      RECT 0.431 0.988 1.265 1.038 ;
      RECT 1.191 1.038 1.241 1.314 ;
      RECT 1.215 0.381 1.265 0.988 ;
      RECT 0.431 0.779 0.521 0.829 ;
      RECT 0.431 0.579 0.521 0.629 ;
      RECT 0.431 1.038 0.481 1.216 ;
      RECT 0.431 0.829 0.481 0.988 ;
      RECT 0.431 0.455 0.481 0.579 ;
      RECT 0.471 0.629 0.521 0.779 ;
      RECT 2.249 0.23 3.141 0.28 ;
      RECT 3.091 0.152 3.141 0.23 ;
      RECT 2.098 0.314 2.299 0.364 ;
      RECT 1.859 0.568 2.148 0.618 ;
      RECT 2.467 0.198 2.549 0.23 ;
      RECT 2.249 0.28 2.299 0.314 ;
      RECT 2.098 0.364 2.148 0.568 ;
      RECT 1.343 0.668 2.245 0.718 ;
      RECT 1.343 0.434 1.561 0.484 ;
      RECT 1.343 1.158 1.713 1.208 ;
      RECT 1.343 0.355 1.393 0.434 ;
      RECT 1.343 1.208 1.393 1.314 ;
      RECT 1.343 0.718 1.393 1.158 ;
      RECT 1.343 0.484 1.393 0.668 ;
      RECT 2.559 0.438 3.901 0.488 ;
      RECT 3.511 0.704 3.901 0.754 ;
      RECT 3.851 0.488 3.901 0.704 ;
      RECT 3.151 1.208 3.561 1.258 ;
      RECT 2.559 0.488 2.609 1.165 ;
      RECT 2.862 0.488 2.912 0.766 ;
      RECT 2.862 0.766 3.005 0.816 ;
      RECT 3.511 0.754 3.561 1.208 ;
      RECT 1.859 0.786 2.381 0.836 ;
      RECT 2.331 0.621 2.381 0.786 ;
      RECT 3.055 0.604 3.765 0.654 ;
      RECT 2.694 0.978 3.105 1.028 ;
      RECT 2.694 0.538 2.801 0.588 ;
      RECT 3.055 0.654 3.105 0.978 ;
      RECT 2.694 0.588 2.744 0.978 ;
      RECT 2.255 1.308 2.457 1.358 ;
      RECT 1.55 1.001 2.497 1.051 ;
      RECT 2.407 0.509 2.497 0.559 ;
      RECT 2.224 0.42 2.457 0.47 ;
      RECT 2.255 1.101 2.305 1.308 ;
      RECT 2.407 1.051 2.457 1.308 ;
      RECT 2.447 0.559 2.497 1.001 ;
      RECT 2.407 0.47 2.457 0.509 ;
      RECT 2.407 0.371 2.457 0.42 ;
      RECT 1.419 1.478 1.941 1.528 ;
      RECT 1.419 1.528 1.469 1.565 ;
      RECT 1.087 1.526 1.317 1.576 ;
      RECT 2.027 1.428 2.077 1.554 ;
      RECT 1.267 1.428 1.317 1.526 ;
      RECT 1.267 1.378 2.077 1.428 ;
      RECT 0.583 0.618 1.029 0.668 ;
      RECT 0.583 0.668 0.633 0.914 ;
      RECT 0.583 0.422 0.633 0.618 ;
      RECT 1.039 0.518 1.165 0.568 ;
      RECT 1.039 0.768 1.089 0.914 ;
      RECT 1.039 0.718 1.165 0.768 ;
      RECT 1.039 0.394 1.089 0.518 ;
      RECT 1.115 0.568 1.165 0.718 ;
      RECT 3.074 1.429 3.461 1.479 ;
      RECT 3.238 0.709 3.461 0.759 ;
      RECT 3.238 0.759 3.288 1.099 ;
      RECT 2.683 1.099 3.288 1.149 ;
      RECT 2.507 1.272 2.733 1.322 ;
      RECT 2.315 1.528 2.557 1.578 ;
      RECT 2.507 1.322 2.557 1.528 ;
      RECT 2.683 1.149 2.733 1.272 ;
      RECT 1.479 1.278 1.865 1.328 ;
      RECT 0.781 0.096 1.491 0.146 ;
    LAYER PO ;
      RECT 2.493 0.068 2.523 0.663 ;
      RECT 3.253 0.068 3.283 1.606 ;
      RECT 0.061 0.066 0.091 1.606 ;
      RECT 0.365 0.068 0.395 1.606 ;
      RECT 0.213 0.066 0.243 1.606 ;
      RECT 1.885 0.758 1.915 1.606 ;
      RECT 1.125 0.068 1.155 1.606 ;
      RECT 3.557 0.068 3.587 1.606 ;
      RECT 4.013 0.068 4.043 1.606 ;
      RECT 2.949 0.068 2.979 1.606 ;
      RECT 2.037 0.068 2.067 1.606 ;
      RECT 0.669 0.068 0.699 1.606 ;
      RECT 1.733 0.068 1.763 1.606 ;
      RECT 0.821 0.068 0.851 1.606 ;
      RECT 2.645 0.068 2.675 1.606 ;
      RECT 2.341 0.068 2.371 1.606 ;
      RECT 3.101 0.068 3.131 1.606 ;
      RECT 3.861 0.068 3.891 1.606 ;
      RECT 1.429 0.068 1.459 1.606 ;
      RECT 2.797 0.068 2.827 1.606 ;
      RECT 0.973 0.068 1.003 1.606 ;
      RECT 3.709 0.068 3.739 1.606 ;
      RECT 1.581 0.068 1.611 1.606 ;
      RECT 0.517 0.068 0.547 1.606 ;
      RECT 1.277 0.068 1.307 0.542 ;
      RECT 4.165 0.068 4.195 1.606 ;
      RECT 1.277 0.99 1.307 1.606 ;
      RECT 3.405 1.012 3.435 1.606 ;
      RECT 2.189 0.068 2.219 1.606 ;
      RECT 1.885 0.068 1.915 0.626 ;
      RECT 3.405 0.068 3.435 0.787 ;
      RECT 2.493 0.882 2.523 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 4.371 1.773 ;
  END
END DFFARX1_RVT

MACRO DFFSSRX1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 4.256 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.881 0.857 0.923 ;
      LAYER M1 ;
        RECT 0.795 0.857 0.967 0.977 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 ;
  END D
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.207 0.705 0.249 0.747 ;
      LAYER M1 ;
        RECT 0.097 0.751 0.207 0.825 ;
        RECT 0.097 0.701 0.269 0.751 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 ;
  END SETB
  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.205 0.401 0.247 ;
        RECT 0.511 0.205 0.553 0.247 ;
      LAYER M1 ;
        RECT 0.249 0.201 0.573 0.251 ;
        RECT 0.249 0.097 0.359 0.201 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 ;
  END RSTB
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.119 1.532 1.161 1.574 ;
      LAYER M1 ;
        RECT 1.009 1.465 1.181 1.576 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.931 0.156 3.973 0.198 ;
        RECT 3.931 0.248 3.973 0.29 ;
        RECT 3.931 1.116 3.973 1.158 ;
        RECT 3.931 1.208 3.973 1.25 ;
        RECT 3.931 1.3 3.973 1.342 ;
        RECT 3.931 1.392 3.973 1.434 ;
        RECT 3.931 1.484 3.973 1.526 ;
      LAYER M1 ;
        RECT 3.927 1.119 3.977 1.546 ;
        RECT 3.927 1.069 4.159 1.119 ;
        RECT 4.049 1.009 4.159 1.069 ;
        RECT 4.109 0.31 4.159 1.009 ;
        RECT 3.927 0.26 4.159 0.31 ;
        RECT 3.927 0.136 3.977 0.26 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.627 0.156 3.669 0.198 ;
        RECT 3.627 0.248 3.669 0.29 ;
        RECT 3.627 0.34 3.669 0.382 ;
        RECT 3.627 0.932 3.669 0.974 ;
        RECT 3.627 1.024 3.669 1.066 ;
        RECT 3.627 1.116 3.669 1.158 ;
        RECT 3.627 1.208 3.669 1.25 ;
        RECT 3.627 1.3 3.669 1.342 ;
        RECT 3.627 1.392 3.669 1.434 ;
        RECT 3.627 1.484 3.669 1.526 ;
      LAYER M1 ;
        RECT 3.623 0.858 3.673 1.546 ;
        RECT 3.623 0.808 4.007 0.858 ;
        RECT 3.957 0.511 4.007 0.808 ;
        RECT 3.897 0.427 4.007 0.511 ;
        RECT 3.623 0.377 4.007 0.427 ;
        RECT 3.623 0.136 3.673 0.377 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.131 0.95 0.173 0.992 ;
        RECT 3.779 0.972 3.821 1.014 ;
        RECT 0.435 1 0.477 1.042 ;
        RECT 0.131 1.042 0.173 1.084 ;
        RECT 3.779 1.064 3.821 1.106 ;
        RECT 0.435 1.092 0.477 1.134 ;
        RECT 2.107 1.12 2.149 1.162 ;
        RECT 0.131 1.134 0.173 1.176 ;
        RECT 3.779 1.156 3.821 1.198 ;
        RECT 0.435 1.184 0.477 1.226 ;
        RECT 2.107 1.212 2.149 1.254 ;
        RECT 0.131 1.226 0.173 1.268 ;
        RECT 3.475 1.236 3.517 1.278 ;
        RECT 3.779 1.248 3.821 1.29 ;
        RECT 0.435 1.276 0.477 1.318 ;
        RECT 2.107 1.304 2.149 1.346 ;
        RECT 0.131 1.318 0.173 1.36 ;
        RECT 1.195 1.32 1.237 1.362 ;
        RECT 3.475 1.328 3.517 1.37 ;
        RECT 2.259 1.336 2.301 1.378 ;
        RECT 3.019 1.42 3.061 1.462 ;
        RECT 3.475 1.42 3.517 1.462 ;
        RECT 2.259 1.428 2.301 1.47 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
        RECT 3.095 1.651 3.137 1.693 ;
        RECT 3.247 1.651 3.289 1.693 ;
        RECT 3.399 1.651 3.441 1.693 ;
        RECT 3.551 1.651 3.593 1.693 ;
        RECT 3.703 1.651 3.745 1.693 ;
        RECT 3.855 1.651 3.897 1.693 ;
        RECT 4.007 1.651 4.049 1.693 ;
        RECT 4.159 1.651 4.201 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 4.256 1.702 ;
        RECT 3.511 1.466 3.561 1.642 ;
        RECT 2.999 1.416 3.561 1.466 ;
        RECT 1.253 1.366 1.303 1.642 ;
        RECT 2.255 1.366 2.305 1.642 ;
        RECT 0.127 1.346 0.177 1.642 ;
        RECT 1.153 1.316 1.303 1.366 ;
        RECT 2.103 1.316 2.305 1.366 ;
        RECT 3.775 0.947 3.825 1.642 ;
        RECT 3.471 1.192 3.521 1.416 ;
        RECT 0.127 1.296 0.481 1.346 ;
        RECT 2.103 1.1 2.153 1.316 ;
        RECT 0.127 0.93 0.177 1.296 ;
        RECT 0.431 0.98 0.481 1.296 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 3.399 -0.021 3.441 0.021 ;
        RECT 3.551 -0.021 3.593 0.021 ;
        RECT 3.703 -0.021 3.745 0.021 ;
        RECT 3.855 -0.021 3.897 0.021 ;
        RECT 4.007 -0.021 4.049 0.021 ;
        RECT 4.159 -0.021 4.201 0.021 ;
        RECT 3.779 0.146 3.821 0.188 ;
        RECT 3.019 0.208 3.061 0.25 ;
        RECT 3.779 0.238 3.821 0.28 ;
        RECT 3.475 0.247 3.517 0.289 ;
        RECT 2.107 0.321 2.149 0.363 ;
        RECT 2.259 0.321 2.301 0.363 ;
        RECT 3.475 0.339 3.517 0.381 ;
        RECT 0.131 0.359 0.173 0.401 ;
        RECT 0.435 0.375 0.477 0.417 ;
        RECT 1.195 0.396 1.237 0.438 ;
        RECT 2.107 0.413 2.149 0.455 ;
        RECT 2.259 0.413 2.301 0.455 ;
        RECT 0.131 0.451 0.173 0.493 ;
        RECT 0.435 0.467 0.477 0.509 ;
        RECT 1.195 0.488 1.237 0.53 ;
      LAYER M1 ;
        RECT 0.431 0.405 0.481 0.529 ;
        RECT 0.127 0.405 0.177 0.513 ;
        RECT 0.127 0.355 0.481 0.405 ;
        RECT 1.191 0.351 1.241 0.576 ;
        RECT 2.103 0.351 2.153 0.475 ;
        RECT 2.255 0.351 2.305 0.475 ;
        RECT 1.191 0.301 2.305 0.351 ;
        RECT 2.975 0.204 3.081 0.254 ;
        RECT 3.471 0.03 3.521 0.401 ;
        RECT 0.127 0.03 0.177 0.355 ;
        RECT 3.775 0.03 3.825 0.303 ;
        RECT 1.875 0.03 1.925 0.301 ;
        RECT 2.975 0.03 3.025 0.204 ;
        RECT 0 -0.03 4.256 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.587 1.184 0.629 1.226 ;
      RECT 1.499 0.45 1.541 0.492 ;
      RECT 2.563 1.213 2.605 1.255 ;
      RECT 1.727 1.421 1.769 1.463 ;
      RECT 1.651 1.082 1.693 1.124 ;
      RECT 0.587 1.092 0.629 1.134 ;
      RECT 1.043 0.998 1.085 1.04 ;
      RECT 2.639 1.532 2.681 1.574 ;
      RECT 1.499 1.082 1.541 1.124 ;
      RECT 2.715 1.199 2.757 1.241 ;
      RECT 0.511 0.848 0.553 0.89 ;
      RECT 1.499 0.45 1.541 0.492 ;
      RECT 2.563 0.32 2.605 0.362 ;
      RECT 1.651 0.45 1.693 0.492 ;
      RECT 0.587 1.276 0.629 1.318 ;
      RECT 0.283 1.184 0.325 1.226 ;
      RECT 1.347 0.814 1.389 0.856 ;
      RECT 2.031 1.421 2.073 1.463 ;
      RECT 0.283 1.184 0.325 1.226 ;
      RECT 2.335 0.577 2.377 0.619 ;
      RECT 2.563 1.121 2.605 1.163 ;
      RECT 1.651 0.45 1.693 0.492 ;
      RECT 2.487 1.532 2.529 1.574 ;
      RECT 1.575 1.532 1.617 1.574 ;
      RECT 2.791 1.532 2.833 1.574 ;
      RECT 1.043 0.814 1.085 0.856 ;
      RECT 0.283 0.475 0.325 0.517 ;
      RECT 2.411 0.32 2.453 0.362 ;
      RECT 1.347 0.998 1.389 1.04 ;
      RECT 0.587 0.305 0.629 0.347 ;
      RECT 1.043 0.814 1.085 0.856 ;
      RECT 2.715 0.32 2.757 0.362 ;
      RECT 1.043 0.998 1.085 1.04 ;
      RECT 0.891 0.305 0.933 0.347 ;
      RECT 0.587 1.092 0.629 1.134 ;
      RECT 1.347 0.814 1.389 0.856 ;
      RECT 0.587 1.184 0.629 1.226 ;
      RECT 0.739 0.447 0.781 0.489 ;
      RECT 2.563 1.305 2.605 1.347 ;
      RECT 0.663 0.577 0.705 0.619 ;
      RECT 1.803 1.092 1.845 1.134 ;
      RECT 3.171 0.481 3.213 0.523 ;
      RECT 0.739 1.184 0.781 1.226 ;
      RECT 1.651 0.99 1.693 1.032 ;
      RECT 1.651 0.45 1.693 0.492 ;
      RECT 0.967 0.108 1.009 0.15 ;
      RECT 0.739 1.184 0.781 1.226 ;
      RECT 1.347 0.998 1.389 1.04 ;
      RECT 0.891 1.32 0.933 1.362 ;
      RECT 3.247 0.108 3.289 0.15 ;
      RECT 1.043 0.906 1.085 0.948 ;
      RECT 2.563 0.412 2.605 0.454 ;
      RECT 1.499 0.99 1.541 1.032 ;
      RECT 2.943 0.658 2.985 0.7 ;
      RECT 3.855 0.664 3.897 0.706 ;
      RECT 2.031 0.998 2.073 1.04 ;
      RECT 1.423 0.63 1.465 0.672 ;
      RECT 3.703 0.596 3.745 0.638 ;
      RECT 3.399 1.532 3.441 1.574 ;
      RECT 0.739 1.092 0.781 1.134 ;
      RECT 1.803 1.184 1.845 1.226 ;
      RECT 1.651 1.174 1.693 1.216 ;
      RECT 1.043 0.906 1.085 0.948 ;
      RECT 1.575 0.155 1.617 0.197 ;
      RECT 1.043 0.513 1.085 0.555 ;
      RECT 2.411 0.412 2.453 0.454 ;
      RECT 1.347 0.45 1.389 0.492 ;
      RECT 1.043 0.421 1.085 0.463 ;
      RECT 1.499 0.45 1.541 0.492 ;
      RECT 1.879 0.777 1.921 0.819 ;
      RECT 0.587 1 0.629 1.042 ;
      RECT 3.399 0.681 3.441 0.723 ;
      RECT 0.587 1 0.629 1.042 ;
      RECT 0.967 0.63 1.009 0.672 ;
      RECT 1.347 1.09 1.389 1.132 ;
      RECT 3.247 0.581 3.289 0.623 ;
      RECT 1.727 0.108 1.769 0.15 ;
      RECT 1.803 0.45 1.845 0.492 ;
      RECT 1.499 1.174 1.541 1.216 ;
      RECT 2.031 0.677 2.073 0.719 ;
      RECT 2.867 1.104 2.909 1.146 ;
      RECT 1.271 0.63 1.313 0.672 ;
      RECT 0.359 1.453 0.401 1.495 ;
      RECT 3.095 0.108 3.137 0.15 ;
      RECT 0.283 1 0.325 1.042 ;
      RECT 0.283 1.092 0.325 1.134 ;
      RECT 0.283 1 0.325 1.042 ;
      RECT 2.411 1.104 2.453 1.146 ;
      RECT 1.347 0.45 1.389 0.492 ;
      RECT 2.639 0.155 2.681 0.197 ;
      RECT 3.171 1.22 3.213 1.262 ;
      RECT 2.791 0.108 2.833 0.15 ;
      RECT 1.043 1.09 1.085 1.132 ;
      RECT 0.739 1.092 0.781 1.134 ;
      RECT 1.347 0.45 1.389 0.492 ;
      RECT 2.031 0.155 2.073 0.197 ;
      RECT 1.347 0.906 1.389 0.948 ;
      RECT 0.283 1.092 0.325 1.134 ;
      RECT 1.347 0.906 1.389 0.948 ;
      RECT 2.867 0.308 2.909 0.35 ;
      RECT 1.423 1.532 1.465 1.574 ;
      RECT 2.715 0.412 2.757 0.454 ;
      RECT 0.663 1.453 0.705 1.495 ;
    LAYER M1 ;
      RECT 1.343 0.726 1.445 0.776 ;
      RECT 1.327 0.446 1.445 0.496 ;
      RECT 1.395 0.626 1.485 0.676 ;
      RECT 1.343 0.776 1.393 1.152 ;
      RECT 1.395 0.676 1.445 0.726 ;
      RECT 1.395 0.496 1.445 0.626 ;
      RECT 3.127 0.477 3.749 0.527 ;
      RECT 3.699 0.527 3.749 0.658 ;
      RECT 2.711 1.216 3.257 1.266 ;
      RECT 2.711 0.3 2.761 1.216 ;
      RECT 2.923 0.654 3.177 0.677 ;
      RECT 3.127 0.704 3.257 0.727 ;
      RECT 2.923 0.677 3.257 0.704 ;
      RECT 3.207 0.727 3.257 1.216 ;
      RECT 3.127 0.527 3.177 0.654 ;
      RECT 1.495 0.726 1.585 0.776 ;
      RECT 1.495 0.526 1.585 0.576 ;
      RECT 0.735 1.202 1.545 1.252 ;
      RECT 1.495 0.43 1.545 0.526 ;
      RECT 1.535 0.576 1.585 0.726 ;
      RECT 1.495 0.776 1.545 1.202 ;
      RECT 0.695 0.752 0.854 0.802 ;
      RECT 0.719 0.443 0.854 0.493 ;
      RECT 0.804 0.493 0.854 0.752 ;
      RECT 0.695 0.802 0.745 1.047 ;
      RECT 0.735 1.097 0.785 1.202 ;
      RECT 0.695 1.047 0.785 1.097 ;
      RECT 2.705 0.104 2.853 0.151 ;
      RECT 2.011 0.154 2.755 0.201 ;
      RECT 2.011 0.151 2.853 0.154 ;
      RECT 0.548 0.573 0.725 0.623 ;
      RECT 0.279 0.844 0.598 0.894 ;
      RECT 0.548 0.623 0.598 0.844 ;
      RECT 0.279 0.601 0.369 0.651 ;
      RECT 0.279 0.455 0.329 0.601 ;
      RECT 0.319 0.651 0.369 0.844 ;
      RECT 0.279 0.894 0.329 1.246 ;
      RECT 1.854 0.773 2.609 0.823 ;
      RECT 2.559 0.823 2.609 1.38 ;
      RECT 2.407 0.823 2.457 1.166 ;
      RECT 2.407 0.3 2.457 0.452 ;
      RECT 2.407 0.452 2.609 0.502 ;
      RECT 2.559 0.502 2.609 0.773 ;
      RECT 2.559 0.3 2.609 0.452 ;
      RECT 2.659 1.316 3.421 1.366 ;
      RECT 3.371 0.677 3.461 0.727 ;
      RECT 3.371 0.727 3.421 1.316 ;
      RECT 2.251 1.216 2.465 1.266 ;
      RECT 2.011 0.994 2.301 1.044 ;
      RECT 2.415 1.528 2.709 1.578 ;
      RECT 2.251 1.044 2.301 1.216 ;
      RECT 2.415 1.266 2.465 1.528 ;
      RECT 2.659 1.366 2.709 1.528 ;
      RECT 1.647 0.573 2.397 0.623 ;
      RECT 1.647 1.196 1.849 1.246 ;
      RECT 1.799 1.072 1.849 1.196 ;
      RECT 1.799 0.43 1.849 0.573 ;
      RECT 1.647 0.623 1.697 1.196 ;
      RECT 1.647 0.43 1.697 0.573 ;
      RECT 3.599 0.708 3.901 0.758 ;
      RECT 3.227 0.577 3.649 0.627 ;
      RECT 3.851 0.621 3.901 0.708 ;
      RECT 3.599 0.627 3.649 0.708 ;
      RECT 2.771 1.528 3.461 1.578 ;
      RECT 3.075 0.104 3.309 0.154 ;
      RECT 2.823 0.304 3.226 0.354 ;
      RECT 3.176 0.154 3.226 0.304 ;
      RECT 2.823 0.808 2.913 0.858 ;
      RECT 2.863 0.858 2.913 1.166 ;
      RECT 2.823 0.354 2.873 0.808 ;
      RECT 0.567 0.301 0.953 0.351 ;
      RECT 0.583 1.316 0.954 1.366 ;
      RECT 0.583 0.98 0.633 1.316 ;
      RECT 1.747 0.88 1.949 0.93 ;
      RECT 1.747 0.673 2.093 0.723 ;
      RECT 1.403 1.528 1.657 1.578 ;
      RECT 1.607 1.367 1.657 1.528 ;
      RECT 1.607 1.317 1.949 1.367 ;
      RECT 1.899 0.93 1.949 1.317 ;
      RECT 1.747 0.723 1.797 0.88 ;
      RECT 0.947 0.104 1.789 0.154 ;
      RECT 1.571 0.154 1.621 0.217 ;
      RECT 0.947 0.626 1.333 0.676 ;
      RECT 1.039 0.676 1.089 1.152 ;
      RECT 1.039 0.401 1.089 0.626 ;
      RECT 1.707 1.417 2.093 1.467 ;
      RECT 0.339 1.449 0.725 1.499 ;
    LAYER PO ;
      RECT 0.669 0.076 0.699 0.651 ;
      RECT 1.581 0.92 1.611 1.606 ;
      RECT 1.429 0.076 1.459 1.606 ;
      RECT 1.885 0.076 1.915 1.606 ;
      RECT 3.709 0.076 3.739 1.606 ;
      RECT 1.277 0.076 1.307 1.606 ;
      RECT 2.341 0.076 2.371 1.606 ;
      RECT 3.405 1.132 3.435 1.606 ;
      RECT 2.037 0.076 2.067 0.751 ;
      RECT 2.949 0.076 2.979 1.606 ;
      RECT 3.253 0.076 3.283 1.606 ;
      RECT 1.733 0.076 1.763 1.606 ;
      RECT 3.861 0.076 3.891 1.606 ;
      RECT 3.101 0.076 3.131 1.606 ;
      RECT 0.973 0.076 1.003 1.606 ;
      RECT 2.645 0.076 2.675 0.597 ;
      RECT 2.493 0.076 2.523 1.606 ;
      RECT 0.517 0.076 0.547 0.597 ;
      RECT 0.517 0.816 0.547 1.606 ;
      RECT 2.797 0.076 2.827 1.606 ;
      RECT 0.821 0.076 0.851 1.606 ;
      RECT 0.061 0.076 0.091 1.606 ;
      RECT 0.213 0.076 0.243 1.606 ;
      RECT 2.037 0.966 2.067 1.606 ;
      RECT 1.125 0.076 1.155 1.606 ;
      RECT 4.165 0.076 4.195 1.606 ;
      RECT 2.189 0.076 2.219 1.606 ;
      RECT 0.669 0.87 0.699 1.606 ;
      RECT 1.581 0.076 1.611 0.597 ;
      RECT 2.645 1.032 2.675 1.606 ;
      RECT 4.013 0.076 4.043 1.606 ;
      RECT 0.365 0.076 0.395 1.606 ;
      RECT 3.405 0.076 3.435 0.755 ;
      RECT 3.557 0.076 3.587 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 4.371 1.773 ;
  END
END DFFSSRX1_RVT

MACRO DFFASX1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 4.256 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.684 0.401 0.726 ;
      LAYER M1 ;
        RECT 0.249 0.68 0.421 0.73 ;
        RECT 0.249 0.553 0.359 0.68 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 ;
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 1.53 0.705 1.572 ;
      LAYER M1 ;
        RECT 0.553 1.424 0.725 1.576 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.247 0.99 3.289 1.032 ;
      LAYER M1 ;
        RECT 3.227 0.857 3.399 1.034 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0441 ;
  END SETB
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.627 0.195 3.669 0.237 ;
        RECT 3.627 0.287 3.669 0.329 ;
        RECT 3.627 0.932 3.669 0.974 ;
        RECT 3.627 1.024 3.669 1.066 ;
        RECT 3.627 1.116 3.669 1.158 ;
        RECT 3.627 1.208 3.669 1.25 ;
        RECT 3.627 1.3 3.669 1.342 ;
        RECT 3.627 1.392 3.669 1.434 ;
        RECT 3.627 1.484 3.669 1.526 ;
      LAYER M1 ;
        RECT 3.897 1.009 4.007 1.119 ;
        RECT 3.623 0.854 3.673 1.546 ;
        RECT 3.957 0.854 4.007 1.009 ;
        RECT 3.623 0.804 4.007 0.854 ;
        RECT 3.957 0.359 4.007 0.804 ;
        RECT 3.623 0.309 4.007 0.359 ;
        RECT 3.623 0.148 3.673 0.309 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.931 0.158 3.973 0.2 ;
        RECT 3.931 1.3 3.973 1.342 ;
        RECT 3.931 1.392 3.973 1.434 ;
        RECT 3.931 1.484 3.973 1.526 ;
      LAYER M1 ;
        RECT 3.927 1.271 3.977 1.546 ;
        RECT 3.927 1.221 4.16 1.271 ;
        RECT 4.05 1.161 4.16 1.221 ;
        RECT 4.109 0.204 4.159 1.161 ;
        RECT 3.911 0.154 4.159 0.204 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.062 0.325 1.104 ;
        RECT 3.779 1.072 3.821 1.114 ;
        RECT 0.739 1.108 0.781 1.15 ;
        RECT 0.891 1.122 0.933 1.164 ;
        RECT 0.283 1.154 0.325 1.196 ;
        RECT 3.779 1.164 3.821 1.206 ;
        RECT 0.739 1.2 0.781 1.242 ;
        RECT 0.891 1.214 0.933 1.256 ;
        RECT 3.779 1.256 3.821 1.298 ;
        RECT 1.803 1.273 1.845 1.315 ;
        RECT 2.107 1.275 2.149 1.317 ;
        RECT 0.739 1.292 0.781 1.334 ;
        RECT 0.891 1.306 0.933 1.348 ;
        RECT 2.867 1.312 2.909 1.354 ;
        RECT 3.475 1.312 3.517 1.354 ;
        RECT 3.779 1.348 3.821 1.39 ;
        RECT 0.891 1.398 0.933 1.44 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
        RECT 3.095 1.651 3.137 1.693 ;
        RECT 3.247 1.651 3.289 1.693 ;
        RECT 3.399 1.651 3.441 1.693 ;
        RECT 3.551 1.651 3.593 1.693 ;
        RECT 3.703 1.651 3.745 1.693 ;
        RECT 3.855 1.651 3.897 1.693 ;
        RECT 4.007 1.651 4.049 1.693 ;
        RECT 4.159 1.651 4.201 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 4.256 1.702 ;
        RECT 3.511 1.358 3.561 1.642 ;
        RECT 0.887 1.354 0.937 1.642 ;
        RECT 1.975 1.321 2.025 1.642 ;
        RECT 2.834 1.308 3.561 1.358 ;
        RECT 0.279 1.033 0.329 1.642 ;
        RECT 3.775 0.947 3.825 1.642 ;
        RECT 0.735 1.304 0.937 1.354 ;
        RECT 1.774 1.271 2.184 1.321 ;
        RECT 0.735 1.088 0.785 1.304 ;
        RECT 0.887 1.101 0.937 1.304 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 3.399 -0.021 3.441 0.021 ;
        RECT 3.551 -0.021 3.593 0.021 ;
        RECT 3.703 -0.021 3.745 0.021 ;
        RECT 3.855 -0.021 3.897 0.021 ;
        RECT 4.007 -0.021 4.049 0.021 ;
        RECT 4.159 -0.021 4.201 0.021 ;
        RECT 3.779 0.158 3.821 0.2 ;
        RECT 0.739 0.2 0.781 0.242 ;
        RECT 1.803 0.217 1.845 0.259 ;
        RECT 0.891 0.275 0.933 0.317 ;
        RECT 1.955 0.307 1.997 0.349 ;
        RECT 1.803 0.309 1.845 0.351 ;
        RECT 0.283 0.344 0.325 0.386 ;
        RECT 2.867 0.347 2.909 0.389 ;
        RECT 3.475 0.347 3.517 0.389 ;
        RECT 0.739 0.388 0.781 0.43 ;
        RECT 0.891 0.388 0.933 0.43 ;
        RECT 1.955 0.399 1.997 0.441 ;
      LAYER M1 ;
        RECT 2.845 0.343 3.537 0.393 ;
        RECT 0.735 0.246 0.785 0.45 ;
        RECT 0.887 0.246 0.937 0.45 ;
        RECT 0.586 0.196 0.937 0.246 ;
        RECT 1.951 0.03 2.001 0.461 ;
        RECT 0.279 0.03 0.329 0.419 ;
        RECT 1.799 0.03 1.849 0.371 ;
        RECT 3.471 0.03 3.521 0.343 ;
        RECT 3.775 0.03 3.825 0.22 ;
        RECT 0.586 0.03 0.636 0.196 ;
        RECT 0 -0.03 4.256 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 2.715 0.547 2.757 0.589 ;
      RECT 1.423 0.098 1.465 0.14 ;
      RECT 1.043 0.852 1.085 0.894 ;
      RECT 2.411 0.391 2.453 0.433 ;
      RECT 3.703 0.608 3.745 0.65 ;
      RECT 1.955 1.17 1.997 1.212 ;
      RECT 1.043 0.76 1.085 0.802 ;
      RECT 0.815 0.622 0.857 0.664 ;
      RECT 2.411 1.291 2.453 1.333 ;
      RECT 0.435 1.154 0.477 1.196 ;
      RECT 2.563 1.103 2.605 1.145 ;
      RECT 2.259 0.391 2.301 0.433 ;
      RECT 0.967 0.622 1.009 0.664 ;
      RECT 3.247 1.415 3.289 1.457 ;
      RECT 1.195 0.319 1.237 0.361 ;
      RECT 2.183 1.532 2.225 1.574 ;
      RECT 2.411 1.199 2.453 1.241 ;
      RECT 3.019 1.212 3.061 1.254 ;
      RECT 2.715 0.979 2.757 1.021 ;
      RECT 0.587 0.442 0.629 0.484 ;
      RECT 0.587 0.442 0.629 0.484 ;
      RECT 1.271 0.1 1.313 0.142 ;
      RECT 0.587 0.442 0.629 0.484 ;
      RECT 1.347 0.375 1.389 0.417 ;
      RECT 1.347 0.375 1.389 0.417 ;
      RECT 1.195 0.319 1.237 0.361 ;
      RECT 1.195 0.319 1.237 0.361 ;
      RECT 0.587 0.852 0.629 0.894 ;
      RECT 3.399 0.713 3.441 0.755 ;
      RECT 1.727 0.542 1.769 0.584 ;
      RECT 0.435 1.154 0.477 1.196 ;
      RECT 0.435 1.062 0.477 1.104 ;
      RECT 1.347 0.375 1.389 0.417 ;
      RECT 1.195 1.252 1.237 1.294 ;
      RECT 1.043 0.506 1.085 0.548 ;
      RECT 0.435 1.062 0.477 1.104 ;
      RECT 1.043 0.414 1.085 0.456 ;
      RECT 2.259 1.199 2.301 1.241 ;
      RECT 3.323 1.212 3.365 1.254 ;
      RECT 2.259 1.291 2.301 1.333 ;
      RECT 3.171 1.112 3.213 1.154 ;
      RECT 1.499 1.16 1.541 1.202 ;
      RECT 1.347 1.16 1.389 1.202 ;
      RECT 1.119 1.53 1.161 1.572 ;
      RECT 0.587 0.76 0.629 0.802 ;
      RECT 2.031 0.644 2.073 0.686 ;
      RECT 2.411 1.107 2.453 1.149 ;
      RECT 3.399 1.538 3.441 1.58 ;
      RECT 2.335 1.432 2.377 1.474 ;
      RECT 1.271 1.49 1.313 1.532 ;
      RECT 2.943 1.538 2.985 1.58 ;
      RECT 3.855 0.608 3.897 0.65 ;
      RECT 3.019 0.447 3.061 0.489 ;
      RECT 2.563 0.49 2.605 0.532 ;
      RECT 2.335 0.76 2.377 0.802 ;
      RECT 2.943 0.188 2.985 0.23 ;
      RECT 2.487 0.18 2.529 0.222 ;
      RECT 1.423 1.501 1.465 1.543 ;
      RECT 3.095 0.608 3.137 0.65 ;
      RECT 1.879 1.478 1.921 1.52 ;
      RECT 1.575 1.003 1.617 1.045 ;
      RECT 1.879 0.542 1.921 0.584 ;
      RECT 1.727 0.76 1.769 0.802 ;
      RECT 2.791 0.647 2.833 0.689 ;
      RECT 1.727 1.48 1.769 1.522 ;
      RECT 1.499 0.436 1.541 0.478 ;
      RECT 0.815 0.1 0.857 0.142 ;
      RECT 1.119 0.649 1.161 0.691 ;
      RECT 0.435 0.492 0.477 0.534 ;
      RECT 1.195 1.16 1.237 1.202 ;
      RECT 2.487 1.432 2.529 1.474 ;
      RECT 1.347 1.252 1.389 1.294 ;
    LAYER M1 ;
      RECT 1.191 0.299 1.281 0.381 ;
      RECT 0.431 0.988 1.265 1.038 ;
      RECT 1.191 1.038 1.241 1.314 ;
      RECT 1.215 0.381 1.265 0.988 ;
      RECT 0.431 0.779 0.521 0.829 ;
      RECT 0.431 0.579 0.521 0.629 ;
      RECT 0.431 1.038 0.481 1.216 ;
      RECT 0.431 0.829 0.481 0.988 ;
      RECT 0.431 0.455 0.481 0.579 ;
      RECT 0.471 0.629 0.521 0.779 ;
      RECT 2.143 0.23 2.989 0.28 ;
      RECT 2.939 0.166 2.989 0.23 ;
      RECT 1.706 0.538 2.193 0.588 ;
      RECT 2.467 0.178 2.549 0.23 ;
      RECT 2.143 0.588 2.193 0.59 ;
      RECT 2.143 0.28 2.193 0.538 ;
      RECT 1.698 0.756 2.397 0.806 ;
      RECT 3.511 0.704 3.901 0.754 ;
      RECT 2.559 0.443 3.901 0.493 ;
      RECT 3.851 0.493 3.901 0.704 ;
      RECT 3.851 0.438 3.901 0.443 ;
      RECT 3.151 1.108 3.561 1.158 ;
      RECT 3.511 0.754 3.561 1.108 ;
      RECT 2.559 0.643 2.853 0.693 ;
      RECT 2.559 0.693 2.609 1.165 ;
      RECT 2.559 0.493 2.609 0.643 ;
      RECT 2.559 0.438 2.609 0.443 ;
      RECT 1.343 0.64 2.093 0.69 ;
      RECT 1.343 0.432 1.561 0.482 ;
      RECT 1.343 1.156 1.561 1.206 ;
      RECT 1.343 0.355 1.393 0.432 ;
      RECT 1.343 0.482 1.393 0.64 ;
      RECT 1.343 1.206 1.393 1.314 ;
      RECT 1.343 0.69 1.393 1.156 ;
      RECT 2.932 0.604 3.765 0.654 ;
      RECT 2.688 0.975 2.982 1.025 ;
      RECT 2.932 0.654 2.982 0.975 ;
      RECT 2.932 0.593 2.982 0.604 ;
      RECT 2.695 0.543 2.982 0.593 ;
      RECT 1.55 1.001 2.497 1.051 ;
      RECT 2.407 0.606 2.497 0.656 ;
      RECT 2.255 1.308 2.457 1.358 ;
      RECT 1.934 1.166 2.305 1.216 ;
      RECT 2.447 0.656 2.497 1.001 ;
      RECT 2.255 0.371 2.305 0.446 ;
      RECT 2.255 0.446 2.457 0.496 ;
      RECT 2.407 1.051 2.457 1.308 ;
      RECT 2.255 1.216 2.305 1.308 ;
      RECT 2.407 0.496 2.457 0.606 ;
      RECT 2.407 0.371 2.457 0.446 ;
      RECT 1.419 1.476 1.789 1.526 ;
      RECT 1.419 1.526 1.469 1.563 ;
      RECT 1.099 1.526 1.317 1.576 ;
      RECT 1.875 1.426 1.925 1.54 ;
      RECT 1.267 1.376 1.925 1.426 ;
      RECT 1.267 1.426 1.317 1.526 ;
      RECT 2.922 1.534 3.461 1.584 ;
      RECT 0.583 0.618 1.029 0.668 ;
      RECT 0.583 0.668 0.633 0.914 ;
      RECT 0.583 0.422 0.633 0.618 ;
      RECT 1.039 0.518 1.165 0.568 ;
      RECT 1.039 0.768 1.089 0.914 ;
      RECT 1.039 0.718 1.165 0.768 ;
      RECT 1.039 0.394 1.089 0.518 ;
      RECT 1.115 0.568 1.165 0.718 ;
      RECT 2.134 1.528 2.682 1.578 ;
      RECT 2.632 1.461 2.682 1.528 ;
      RECT 2.632 1.411 3.309 1.461 ;
      RECT 3.051 0.709 3.461 0.759 ;
      RECT 3.051 0.759 3.101 1.099 ;
      RECT 2.683 1.099 3.101 1.149 ;
      RECT 2.507 1.272 2.733 1.322 ;
      RECT 2.315 1.428 2.557 1.478 ;
      RECT 2.507 1.322 2.557 1.428 ;
      RECT 2.683 1.149 2.733 1.272 ;
      RECT 2.683 1.096 2.733 1.099 ;
      RECT 0.795 0.096 1.491 0.146 ;
      RECT 2.999 1.208 3.385 1.258 ;
    LAYER PO ;
      RECT 3.405 1.012 3.435 1.606 ;
      RECT 2.493 0.068 2.523 0.622 ;
      RECT 0.061 0.066 0.091 1.606 ;
      RECT 0.365 0.068 0.395 1.606 ;
      RECT 0.213 0.066 0.243 1.606 ;
      RECT 1.125 0.068 1.155 1.606 ;
      RECT 3.557 0.068 3.587 1.606 ;
      RECT 4.013 0.068 4.043 1.606 ;
      RECT 2.189 0.068 2.219 1.606 ;
      RECT 3.253 0.068 3.283 1.606 ;
      RECT 0.669 0.068 0.699 1.606 ;
      RECT 2.037 0.068 2.067 1.606 ;
      RECT 0.821 0.068 0.851 1.606 ;
      RECT 2.645 0.068 2.675 1.606 ;
      RECT 2.341 0.068 2.371 1.606 ;
      RECT 2.949 0.068 2.979 1.606 ;
      RECT 3.861 0.068 3.891 1.606 ;
      RECT 3.101 0.068 3.131 1.606 ;
      RECT 0.973 0.068 1.003 1.606 ;
      RECT 3.709 0.068 3.739 1.606 ;
      RECT 0.517 0.068 0.547 1.606 ;
      RECT 1.277 0.068 1.307 0.542 ;
      RECT 4.165 0.068 4.195 1.606 ;
      RECT 1.277 0.99 1.307 1.606 ;
      RECT 1.733 0.728 1.763 1.604 ;
      RECT 1.885 0.066 1.915 1.604 ;
      RECT 3.405 0.068 3.435 0.787 ;
      RECT 2.797 0.065 2.827 1.603 ;
      RECT 1.581 0.066 1.611 1.604 ;
      RECT 1.429 0.066 1.459 1.604 ;
      RECT 1.733 0.066 1.763 0.616 ;
      RECT 2.493 0.882 2.523 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 4.371 1.773 ;
      RECT 2.66 0.669 2.964 0.679 ;
  END
END DFFASX1_RVT

MACRO NAND2X0_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.912 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.043 0.553 1.085 ;
      LAYER M1 ;
        RECT 0.401 1.089 0.506 1.119 ;
        RECT 0.401 1.039 0.573 1.089 ;
        RECT 0.401 1.009 0.506 1.039 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0186 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.254 0.785 0.359 0.815 ;
        RECT 0.254 0.735 0.426 0.785 ;
        RECT 0.254 0.705 0.359 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0186 ;
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.587 0.141 0.629 0.183 ;
        RECT 0.587 0.233 0.629 0.275 ;
        RECT 0.587 0.325 0.629 0.367 ;
        RECT 0.283 1.305 0.325 1.347 ;
        RECT 0.587 1.305 0.629 1.347 ;
        RECT 0.283 1.397 0.325 1.439 ;
        RECT 0.587 1.397 0.629 1.439 ;
        RECT 0.283 1.489 0.325 1.531 ;
        RECT 0.587 1.489 0.629 1.531 ;
      LAYER M1 ;
        RECT 0.279 1.235 0.329 1.551 ;
        RECT 0.583 1.235 0.633 1.551 ;
        RECT 0.279 1.185 0.673 1.235 ;
        RECT 0.623 0.967 0.673 1.185 ;
        RECT 0.553 0.857 0.673 0.967 ;
        RECT 0.623 0.671 0.673 0.857 ;
        RECT 0.583 0.621 0.673 0.671 ;
        RECT 0.583 0.106 0.633 0.621 ;
    END
    ANTENNADIFFAREA 0.0938 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.435 1.305 0.477 1.347 ;
        RECT 0.435 1.397 0.477 1.439 ;
        RECT 0.435 1.489 0.477 1.531 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 0.912 1.702 ;
        RECT 0.431 1.285 0.481 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.283 0.141 0.325 0.183 ;
        RECT 0.283 0.233 0.325 0.275 ;
        RECT 0.283 0.325 0.325 0.367 ;
      LAYER M1 ;
        RECT 0.279 0.03 0.329 0.402 ;
        RECT 0 -0.03 0.912 0.03 ;
    END
  END VSS
  OBS
    LAYER PO ;
      RECT 0.669 0.071 0.699 1.601 ;
      RECT 0.365 0.071 0.395 1.601 ;
      RECT 0.517 0.071 0.547 1.601 ;
      RECT 0.213 0.071 0.243 1.601 ;
      RECT 0.821 0.071 0.851 1.601 ;
      RECT 0.061 0.071 0.091 1.601 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.027 1.773 ;
  END
END NAND2X0_RVT

MACRO AO21X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.89 0.553 0.932 ;
      LAYER M1 ;
        RECT 0.492 0.857 0.663 0.967 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0243 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.725 0.401 0.767 ;
      LAYER M1 ;
        RECT 0.249 0.705 0.421 0.815 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0243 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.117 0.857 0.159 ;
      LAYER M1 ;
        RECT 0.705 0.097 0.877 0.207 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0225 ;
  END A3
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.195 0.154 1.237 0.196 ;
        RECT 1.195 0.246 1.237 0.288 ;
        RECT 1.195 0.338 1.237 0.38 ;
        RECT 1.195 0.43 1.237 0.472 ;
        RECT 1.195 0.848 1.237 0.89 ;
        RECT 1.195 0.94 1.237 0.982 ;
        RECT 1.195 1.032 1.237 1.074 ;
        RECT 1.195 1.124 1.237 1.166 ;
        RECT 1.195 1.216 1.237 1.258 ;
        RECT 1.195 1.308 1.237 1.35 ;
        RECT 1.195 1.4 1.237 1.442 ;
        RECT 1.195 1.492 1.237 1.534 ;
      LAYER M1 ;
        RECT 1.191 1.271 1.241 1.554 ;
        RECT 1.161 1.161 1.271 1.271 ;
        RECT 1.191 0.855 1.241 1.161 ;
        RECT 1.191 0.805 1.281 0.855 ;
        RECT 1.231 0.492 1.281 0.805 ;
        RECT 1.191 0.442 1.281 0.492 ;
        RECT 1.191 0.134 1.241 0.442 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.043 0.848 1.085 0.89 ;
        RECT 1.043 0.94 1.085 0.982 ;
        RECT 1.043 1.032 1.085 1.074 ;
        RECT 1.043 1.124 1.085 1.166 ;
        RECT 0.283 1.133 0.325 1.175 ;
        RECT 1.043 1.216 1.085 1.258 ;
        RECT 0.283 1.225 0.325 1.267 ;
        RECT 0.587 1.225 0.629 1.267 ;
        RECT 1.043 1.308 1.085 1.35 ;
        RECT 0.283 1.317 0.325 1.359 ;
        RECT 0.587 1.317 0.629 1.359 ;
        RECT 1.043 1.4 1.085 1.442 ;
        RECT 0.283 1.409 0.325 1.451 ;
        RECT 0.587 1.409 0.629 1.451 ;
        RECT 1.043 1.492 1.085 1.534 ;
        RECT 0.283 1.501 0.325 1.543 ;
        RECT 0.587 1.501 0.629 1.543 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.52 1.702 ;
        RECT 0.279 1.113 0.329 1.642 ;
        RECT 0.582 1.205 0.632 1.642 ;
        RECT 1.039 0.828 1.089 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.043 0.134 1.085 0.176 ;
        RECT 1.043 0.226 1.085 0.268 ;
        RECT 1.043 0.318 1.085 0.36 ;
        RECT 0.283 0.408 0.325 0.45 ;
        RECT 0.739 0.408 0.781 0.45 ;
        RECT 1.043 0.41 1.085 0.452 ;
        RECT 0.283 0.5 0.325 0.542 ;
        RECT 0.739 0.5 0.781 0.542 ;
      LAYER M1 ;
        RECT 0.279 0.338 0.329 0.562 ;
        RECT 0.735 0.338 0.785 0.562 ;
        RECT 0.279 0.288 0.785 0.338 ;
        RECT 1.04 0.03 1.09 0.472 ;
        RECT 0.279 0.03 0.329 0.288 ;
        RECT 0 -0.03 1.52 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.583 0.62 1.181 0.67 ;
      RECT 0.583 0.388 0.633 0.62 ;
      RECT 0.887 0.67 0.937 1.568 ;
      RECT 0.887 0.388 0.937 0.62 ;
      RECT 0.735 1.12 0.785 1.563 ;
      RECT 0.431 1.07 0.785 1.12 ;
      RECT 0.431 1.12 0.481 1.568 ;
    LAYER PO ;
      RECT 1.277 0.063 1.307 1.604 ;
      RECT 0.213 0.064 0.243 1.613 ;
      RECT 1.125 0.064 1.155 1.604 ;
      RECT 0.821 0.059 0.851 1.613 ;
      RECT 0.973 0.064 1.003 1.613 ;
      RECT 0.669 0.064 0.699 1.613 ;
      RECT 0.061 0.064 0.091 1.613 ;
      RECT 1.429 0.063 1.459 1.604 ;
      RECT 0.365 0.059 0.395 1.613 ;
      RECT 0.517 0.064 0.547 1.613 ;
    LAYER CO ;
      RECT 0.891 1.041 0.933 1.083 ;
      RECT 1.119 0.624 1.161 0.666 ;
      RECT 0.739 1.133 0.781 1.175 ;
      RECT 0.739 1.501 0.781 1.543 ;
      RECT 0.891 1.225 0.933 1.267 ;
      RECT 0.435 1.317 0.477 1.359 ;
      RECT 0.435 1.409 0.477 1.451 ;
      RECT 0.435 1.501 0.477 1.543 ;
      RECT 0.891 0.408 0.933 0.45 ;
      RECT 0.891 1.317 0.933 1.359 ;
      RECT 0.435 1.225 0.477 1.267 ;
      RECT 0.891 1.133 0.933 1.175 ;
      RECT 0.739 1.225 0.781 1.267 ;
      RECT 0.587 0.5 0.629 0.542 ;
      RECT 0.891 1.409 0.933 1.451 ;
      RECT 0.891 1.501 0.933 1.543 ;
      RECT 0.739 1.317 0.781 1.359 ;
      RECT 0.891 0.5 0.933 0.542 ;
      RECT 0.587 0.408 0.629 0.45 ;
      RECT 0.739 1.409 0.781 1.451 ;
      RECT 0.435 1.133 0.477 1.175 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.635 1.773 ;
  END
END AO21X1_RVT

MACRO NAND4X0_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.216 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.891 0.857 0.933 ;
      LAYER M1 ;
        RECT 0.705 0.937 0.815 0.967 ;
        RECT 0.705 0.887 0.877 0.937 ;
        RECT 0.705 0.857 0.815 0.887 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0276 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.738 0.705 0.78 ;
      LAYER M1 ;
        RECT 0.553 0.785 0.663 0.815 ;
        RECT 0.553 0.735 0.725 0.785 ;
        RECT 0.553 0.705 0.663 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0276 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.891 0.553 0.933 ;
      LAYER M1 ;
        RECT 0.401 0.937 0.511 0.967 ;
        RECT 0.401 0.887 0.573 0.937 ;
        RECT 0.401 0.857 0.511 0.887 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0276 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.738 0.401 0.78 ;
      LAYER M1 ;
        RECT 0.249 0.785 0.359 0.815 ;
        RECT 0.249 0.735 0.421 0.785 ;
        RECT 0.249 0.705 0.359 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0276 ;
  END A4
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.891 0.141 0.933 0.183 ;
        RECT 0.891 0.233 0.933 0.275 ;
        RECT 0.891 0.325 0.933 0.367 ;
        RECT 0.891 0.417 0.933 0.459 ;
        RECT 0.891 0.509 0.933 0.551 ;
        RECT 0.283 1.213 0.325 1.255 ;
        RECT 0.587 1.213 0.629 1.255 ;
        RECT 0.891 1.213 0.933 1.255 ;
        RECT 0.283 1.305 0.325 1.347 ;
        RECT 0.587 1.305 0.629 1.347 ;
        RECT 0.891 1.305 0.933 1.347 ;
        RECT 0.283 1.397 0.325 1.439 ;
        RECT 0.587 1.397 0.629 1.439 ;
        RECT 0.891 1.397 0.933 1.439 ;
        RECT 0.283 1.489 0.325 1.531 ;
        RECT 0.587 1.489 0.629 1.531 ;
        RECT 0.891 1.489 0.933 1.531 ;
      LAYER M1 ;
        RECT 0.279 1.103 0.329 1.551 ;
        RECT 0.583 1.103 0.633 1.551 ;
        RECT 0.887 1.103 0.937 1.551 ;
        RECT 0.279 1.053 0.977 1.103 ;
        RECT 0.927 0.815 0.977 1.053 ;
        RECT 0.857 0.705 0.977 0.815 ;
        RECT 0.927 0.651 0.977 0.705 ;
        RECT 0.887 0.601 0.977 0.651 ;
        RECT 0.887 0.121 0.937 0.601 ;
    END
    ANTENNADIFFAREA 0.1834 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.435 1.213 0.477 1.255 ;
        RECT 0.739 1.213 0.781 1.255 ;
        RECT 0.435 1.305 0.477 1.347 ;
        RECT 0.739 1.305 0.781 1.347 ;
        RECT 0.435 1.397 0.477 1.439 ;
        RECT 0.739 1.397 0.781 1.439 ;
        RECT 0.435 1.489 0.477 1.531 ;
        RECT 0.739 1.489 0.781 1.531 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.216 1.702 ;
        RECT 0.431 1.193 0.481 1.642 ;
        RECT 0.735 1.193 0.785 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 0.283 0.141 0.325 0.183 ;
        RECT 0.283 0.233 0.325 0.275 ;
        RECT 0.283 0.325 0.325 0.367 ;
        RECT 0.283 0.417 0.325 0.459 ;
        RECT 0.283 0.509 0.325 0.551 ;
      LAYER M1 ;
        RECT 0.279 0.03 0.329 0.571 ;
        RECT 0 -0.03 1.216 0.03 ;
    END
  END VSS
  OBS
    LAYER PO ;
      RECT 1.125 0.071 1.155 1.61 ;
      RECT 0.973 0.071 1.003 1.61 ;
      RECT 0.669 0.071 0.699 1.61 ;
      RECT 0.365 0.071 0.395 1.61 ;
      RECT 0.517 0.071 0.547 1.61 ;
      RECT 0.213 0.071 0.243 1.61 ;
      RECT 0.821 0.071 0.851 1.61 ;
      RECT 0.061 0.071 0.091 1.61 ;
    LAYER NWELL ;
      RECT -0.115 0.716 1.331 1.773 ;
      RECT -0.115 0.679 0.191 0.716 ;
      RECT 1.018 0.679 1.331 0.716 ;
  END
END NAND4X0_RVT

MACRO AO22X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.744 0.401 0.786 ;
      LAYER M1 ;
        RECT 0.249 0.705 0.404 0.815 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.969 0.553 1.011 ;
      LAYER M1 ;
        RECT 0.401 1.009 0.557 1.119 ;
        RECT 0.507 0.949 0.557 1.009 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.121 0.857 0.163 ;
      LAYER M1 ;
        RECT 0.705 0.097 0.863 0.207 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.6 0.705 0.642 ;
      LAYER M1 ;
        RECT 0.553 0.553 0.708 0.663 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 ;
  END A4
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.195 0.165 1.237 0.207 ;
        RECT 1.195 0.257 1.237 0.299 ;
        RECT 1.195 0.349 1.237 0.391 ;
        RECT 1.195 0.441 1.237 0.483 ;
        RECT 1.195 0.86 1.237 0.902 ;
        RECT 1.195 0.952 1.237 0.994 ;
        RECT 1.195 1.044 1.237 1.086 ;
        RECT 1.195 1.136 1.237 1.178 ;
        RECT 1.195 1.228 1.237 1.27 ;
        RECT 1.195 1.32 1.237 1.362 ;
        RECT 1.195 1.412 1.237 1.454 ;
        RECT 1.195 1.504 1.237 1.546 ;
      LAYER M1 ;
        RECT 1.191 1.271 1.241 1.566 ;
        RECT 1.161 1.161 1.271 1.271 ;
        RECT 1.191 0.865 1.241 1.161 ;
        RECT 1.191 0.815 1.281 0.865 ;
        RECT 1.231 0.504 1.281 0.815 ;
        RECT 1.191 0.438 1.281 0.504 ;
        RECT 1.191 0.145 1.241 0.438 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.043 0.86 1.085 0.902 ;
        RECT 1.043 0.952 1.085 0.994 ;
        RECT 1.043 1.044 1.085 1.086 ;
        RECT 1.043 1.136 1.085 1.178 ;
        RECT 1.043 1.228 1.085 1.27 ;
        RECT 1.043 1.32 1.085 1.362 ;
        RECT 0.435 1.407 0.477 1.449 ;
        RECT 1.043 1.412 1.085 1.454 ;
        RECT 0.435 1.499 0.477 1.541 ;
        RECT 1.043 1.504 1.085 1.546 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.52 1.702 ;
        RECT 0.431 1.387 0.481 1.642 ;
        RECT 1.039 0.84 1.089 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.043 0.165 1.085 0.207 ;
        RECT 1.043 0.257 1.085 0.299 ;
        RECT 0.587 0.34 0.629 0.382 ;
        RECT 1.043 0.349 1.085 0.391 ;
        RECT 1.043 0.441 1.085 0.483 ;
      LAYER M1 ;
        RECT 1.039 0.03 1.089 0.503 ;
        RECT 0.583 0.03 0.633 0.402 ;
        RECT 0 -0.03 1.52 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.758 0.618 1.181 0.668 ;
      RECT 0.279 0.503 0.329 0.57 ;
      RECT 0.279 0.304 0.329 0.453 ;
      RECT 0.735 0.813 0.808 0.863 ;
      RECT 0.758 0.668 0.808 0.813 ;
      RECT 0.735 0.863 0.785 1.237 ;
      RECT 0.887 0.503 0.937 0.568 ;
      RECT 0.279 0.453 0.937 0.503 ;
      RECT 0.887 0.301 0.937 0.453 ;
      RECT 0.758 0.503 0.808 0.618 ;
      RECT 0.583 1.337 0.633 1.572 ;
      RECT 0.279 1.287 0.937 1.337 ;
      RECT 0.887 1.337 0.937 1.571 ;
      RECT 0.279 1.337 0.329 1.571 ;
    LAYER PO ;
      RECT 1.277 0.075 1.307 1.616 ;
      RECT 0.669 0.072 0.699 1.621 ;
      RECT 0.517 0.072 0.547 1.621 ;
      RECT 0.365 0.067 0.395 1.621 ;
      RECT 1.429 0.075 1.459 1.616 ;
      RECT 0.061 0.072 0.091 1.621 ;
      RECT 0.973 0.076 1.003 1.621 ;
      RECT 1.125 0.076 1.155 1.616 ;
      RECT 0.821 0.072 0.851 1.621 ;
      RECT 0.213 0.072 0.243 1.621 ;
    LAYER CO ;
      RECT 0.283 1.325 0.325 1.367 ;
      RECT 0.891 1.325 0.933 1.367 ;
      RECT 0.283 1.417 0.325 1.459 ;
      RECT 0.283 1.509 0.325 1.551 ;
      RECT 0.739 1.175 0.781 1.217 ;
      RECT 0.739 1.083 0.781 1.125 ;
      RECT 0.587 1.509 0.629 1.551 ;
      RECT 0.587 1.417 0.629 1.459 ;
      RECT 0.283 0.508 0.325 0.55 ;
      RECT 0.891 0.506 0.933 0.548 ;
      RECT 0.891 1.509 0.933 1.551 ;
      RECT 1.119 0.622 1.161 0.664 ;
      RECT 0.891 0.414 0.933 0.456 ;
      RECT 0.891 0.322 0.933 0.364 ;
      RECT 0.283 0.324 0.325 0.366 ;
      RECT 0.283 0.416 0.325 0.458 ;
      RECT 0.587 1.325 0.629 1.367 ;
      RECT 0.891 1.417 0.933 1.459 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.635 1.773 ;
  END
END AO22X1_RVT

MACRO AND2X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.216 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.891 0.553 0.933 ;
      LAYER M1 ;
        RECT 0.401 0.937 0.511 0.967 ;
        RECT 0.401 0.887 0.573 0.937 ;
        RECT 0.401 0.857 0.511 0.887 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0243 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.249 0.785 0.359 0.815 ;
        RECT 0.249 0.735 0.421 0.785 ;
        RECT 0.249 0.705 0.359 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0243 ;
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.891 0.15 0.933 0.192 ;
        RECT 0.891 0.242 0.933 0.284 ;
        RECT 0.891 0.334 0.933 0.376 ;
        RECT 0.891 0.426 0.933 0.468 ;
        RECT 0.891 0.93 0.933 0.972 ;
        RECT 0.891 1.022 0.933 1.064 ;
        RECT 0.891 1.114 0.933 1.156 ;
        RECT 0.891 1.206 0.933 1.248 ;
        RECT 0.891 1.298 0.933 1.34 ;
        RECT 0.891 1.39 0.933 1.432 ;
        RECT 0.891 1.482 0.933 1.524 ;
      LAYER M1 ;
        RECT 0.887 0.909 0.937 1.559 ;
        RECT 0.887 0.859 1.024 0.909 ;
        RECT 0.974 0.663 1.024 0.859 ;
        RECT 0.974 0.602 1.119 0.663 ;
        RECT 0.887 0.553 1.119 0.602 ;
        RECT 0.887 0.552 1.045 0.553 ;
        RECT 0.887 0.117 0.937 0.552 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.739 0.93 0.781 0.972 ;
        RECT 0.739 1.022 0.781 1.064 ;
        RECT 0.739 1.114 0.781 1.156 ;
        RECT 0.739 1.206 0.781 1.248 ;
        RECT 0.739 1.298 0.781 1.34 ;
        RECT 0.739 1.39 0.781 1.432 ;
        RECT 0.435 1.4 0.477 1.442 ;
        RECT 0.739 1.482 0.781 1.524 ;
        RECT 0.435 1.492 0.477 1.534 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.216 1.702 ;
        RECT 0.431 1.363 0.481 1.642 ;
        RECT 0.735 0.893 0.785 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 0.283 0.141 0.325 0.183 ;
        RECT 0.739 0.15 0.781 0.192 ;
        RECT 0.283 0.233 0.325 0.275 ;
        RECT 0.739 0.242 0.781 0.284 ;
        RECT 0.283 0.325 0.325 0.367 ;
        RECT 0.739 0.334 0.781 0.376 ;
        RECT 0.283 0.417 0.325 0.459 ;
        RECT 0.739 0.426 0.781 0.468 ;
      LAYER M1 ;
        RECT 0.735 0.03 0.785 0.503 ;
        RECT 0.279 0.03 0.329 0.479 ;
        RECT 0 -0.03 1.216 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.583 0.656 0.877 0.706 ;
      RECT 0.279 1.094 0.329 1.569 ;
      RECT 0.624 0.656 0.674 1.143 ;
      RECT 0.304 1.094 0.672 1.144 ;
      RECT 0.583 1.119 0.633 1.569 ;
      RECT 0.583 0.106 0.633 0.696 ;
    LAYER PO ;
      RECT 0.365 0.071 0.395 1.604 ;
      RECT 0.517 0.071 0.547 1.604 ;
      RECT 0.213 0.071 0.243 1.604 ;
      RECT 0.061 0.071 0.091 1.604 ;
      RECT 0.973 0.072 1.003 1.604 ;
      RECT 1.125 0.072 1.155 1.604 ;
      RECT 0.821 0.072 0.851 1.606 ;
      RECT 0.669 0.071 0.699 1.604 ;
    LAYER CO ;
      RECT 0.283 1.4 0.325 1.442 ;
      RECT 0.283 1.492 0.325 1.534 ;
      RECT 0.587 1.4 0.629 1.442 ;
      RECT 0.587 1.492 0.629 1.534 ;
      RECT 0.587 0.325 0.629 0.367 ;
      RECT 0.587 0.417 0.629 0.459 ;
      RECT 0.283 1.308 0.325 1.35 ;
      RECT 0.587 0.141 0.629 0.183 ;
      RECT 0.587 0.233 0.629 0.275 ;
      RECT 0.283 1.216 0.325 1.258 ;
      RECT 0.587 1.308 0.629 1.35 ;
      RECT 0.587 1.216 0.629 1.258 ;
      RECT 0.815 0.66 0.857 0.702 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.321 1.773 ;
  END
END AND2X1_RVT

MACRO AND3X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.368 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.742 0.705 0.784 ;
      LAYER M1 ;
        RECT 0.553 0.787 0.663 0.815 ;
        RECT 0.553 0.737 0.725 0.787 ;
        RECT 0.553 0.705 0.663 0.737 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0204 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.045 0.553 1.087 ;
      LAYER M1 ;
        RECT 0.401 1.091 0.511 1.119 ;
        RECT 0.401 1.041 0.573 1.091 ;
        RECT 0.401 1.009 0.511 1.041 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0204 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.742 0.401 0.784 ;
      LAYER M1 ;
        RECT 0.249 0.787 0.359 0.815 ;
        RECT 0.249 0.737 0.421 0.787 ;
        RECT 0.249 0.705 0.359 0.737 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0204 ;
  END A3
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.043 0.141 1.085 0.183 ;
        RECT 1.043 0.233 1.085 0.275 ;
        RECT 1.043 0.325 1.085 0.367 ;
        RECT 1.043 0.417 1.085 0.459 ;
        RECT 1.043 0.838 1.085 0.88 ;
        RECT 1.043 0.93 1.085 0.972 ;
        RECT 1.043 1.022 1.085 1.064 ;
        RECT 1.043 1.114 1.085 1.156 ;
        RECT 1.043 1.206 1.085 1.248 ;
        RECT 1.043 1.298 1.085 1.34 ;
        RECT 1.043 1.39 1.085 1.432 ;
        RECT 1.043 1.482 1.085 1.524 ;
      LAYER M1 ;
        RECT 1.039 0.815 1.089 1.544 ;
        RECT 1.039 0.765 1.271 0.815 ;
        RECT 1.116 0.705 1.271 0.765 ;
        RECT 1.116 0.53 1.166 0.705 ;
        RECT 1.039 0.48 1.166 0.53 ;
        RECT 1.039 0.121 1.089 0.48 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.891 0.838 0.933 0.88 ;
        RECT 0.891 0.93 0.933 0.972 ;
        RECT 0.891 1.022 0.933 1.064 ;
        RECT 0.891 1.114 0.933 1.156 ;
        RECT 0.891 1.206 0.933 1.248 ;
        RECT 0.891 1.298 0.933 1.34 ;
        RECT 0.283 1.307 0.325 1.349 ;
        RECT 0.587 1.307 0.629 1.349 ;
        RECT 0.891 1.39 0.933 1.432 ;
        RECT 0.283 1.399 0.325 1.441 ;
        RECT 0.587 1.399 0.629 1.441 ;
        RECT 0.891 1.482 0.933 1.524 ;
        RECT 0.283 1.491 0.325 1.533 ;
        RECT 0.587 1.491 0.629 1.533 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.368 1.702 ;
        RECT 0.279 1.285 0.329 1.642 ;
        RECT 0.583 1.285 0.633 1.642 ;
        RECT 0.887 0.818 0.937 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 0.283 0.141 0.325 0.183 ;
        RECT 0.891 0.141 0.933 0.183 ;
        RECT 0.283 0.233 0.325 0.275 ;
        RECT 0.891 0.233 0.933 0.275 ;
        RECT 0.283 0.325 0.325 0.367 ;
        RECT 0.891 0.325 0.933 0.367 ;
        RECT 0.283 0.417 0.325 0.459 ;
        RECT 0.891 0.417 0.933 0.459 ;
      LAYER M1 ;
        RECT 0.279 0.03 0.329 0.479 ;
        RECT 0.887 0.03 0.937 0.479 ;
        RECT 0 -0.03 1.368 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.784 0.658 1.048 0.708 ;
      RECT 0.431 1.184 0.481 1.553 ;
      RECT 0.775 0.565 0.825 1.234 ;
      RECT 0.735 0.121 0.785 0.614 ;
      RECT 0.456 1.184 0.809 1.234 ;
      RECT 0.735 1.187 0.785 1.553 ;
      RECT 0.735 0.565 0.808 0.615 ;
    LAYER PO ;
      RECT 1.125 0.072 1.155 1.603 ;
      RECT 1.277 0.072 1.307 1.603 ;
      RECT 0.973 0.071 1.003 1.604 ;
      RECT 0.061 0.071 0.091 1.603 ;
      RECT 0.821 0.071 0.851 1.603 ;
      RECT 0.213 0.071 0.243 1.603 ;
      RECT 0.517 0.071 0.547 1.603 ;
      RECT 0.365 0.071 0.395 1.603 ;
      RECT 0.669 0.071 0.699 1.603 ;
    LAYER CO ;
      RECT 0.967 0.662 1.009 0.704 ;
      RECT 0.739 1.491 0.781 1.533 ;
      RECT 0.739 1.307 0.781 1.349 ;
      RECT 0.739 1.399 0.781 1.441 ;
      RECT 0.739 0.141 0.781 0.183 ;
      RECT 0.739 0.233 0.781 0.275 ;
      RECT 0.739 0.325 0.781 0.367 ;
      RECT 0.739 0.417 0.781 0.459 ;
      RECT 0.435 1.491 0.477 1.533 ;
      RECT 0.435 1.399 0.477 1.441 ;
      RECT 0.435 1.307 0.477 1.349 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.483 1.773 ;
  END
END AND3X1_RVT

MACRO DFFX2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 4.256 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.684 0.401 0.726 ;
      LAYER M1 ;
        RECT 0.249 0.68 0.421 0.73 ;
        RECT 0.249 0.553 0.359 0.68 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 ;
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 1.53 0.705 1.572 ;
      LAYER M1 ;
        RECT 0.553 1.424 0.725 1.576 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.475 0.195 3.517 0.237 ;
        RECT 3.475 0.287 3.517 0.329 ;
        RECT 3.475 0.932 3.517 0.974 ;
        RECT 3.475 1.024 3.517 1.066 ;
        RECT 3.475 1.116 3.517 1.158 ;
        RECT 3.475 1.208 3.517 1.25 ;
        RECT 3.475 1.3 3.517 1.342 ;
        RECT 3.475 1.392 3.517 1.434 ;
        RECT 3.475 1.484 3.517 1.526 ;
      LAYER M1 ;
        RECT 3.471 0.854 3.521 1.546 ;
        RECT 3.471 0.804 4.017 0.854 ;
        RECT 3.967 0.511 4.017 0.804 ;
        RECT 3.897 0.444 4.017 0.511 ;
        RECT 3.471 0.394 4.017 0.444 ;
        RECT 3.471 0.148 3.521 0.394 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.779 0.195 3.821 0.237 ;
        RECT 3.779 1.024 3.821 1.066 ;
        RECT 3.779 1.116 3.821 1.158 ;
        RECT 3.779 1.208 3.821 1.25 ;
        RECT 3.779 1.3 3.821 1.342 ;
        RECT 3.779 1.392 3.821 1.434 ;
        RECT 3.779 1.484 3.821 1.526 ;
      LAYER M1 ;
        RECT 3.775 0.968 3.825 1.546 ;
        RECT 3.775 0.918 4.141 0.968 ;
        RECT 4.091 0.32 4.141 0.918 ;
        RECT 3.775 0.27 4.141 0.32 ;
        RECT 3.775 0.148 3.825 0.27 ;
        RECT 4.091 0.207 4.141 0.27 ;
        RECT 4.049 0.097 4.159 0.207 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 3.323 0.932 3.365 0.974 ;
        RECT 3.627 0.98 3.669 1.022 ;
        RECT 3.323 1.024 3.365 1.066 ;
        RECT 0.283 1.062 0.325 1.104 ;
        RECT 3.627 1.072 3.669 1.114 ;
        RECT 3.931 1.072 3.973 1.114 ;
        RECT 0.739 1.108 0.781 1.15 ;
        RECT 3.323 1.116 3.365 1.158 ;
        RECT 0.891 1.122 0.933 1.164 ;
        RECT 0.283 1.154 0.325 1.196 ;
        RECT 3.627 1.164 3.669 1.206 ;
        RECT 3.931 1.164 3.973 1.206 ;
        RECT 0.739 1.2 0.781 1.242 ;
        RECT 3.323 1.208 3.365 1.25 ;
        RECT 0.891 1.214 0.933 1.256 ;
        RECT 3.627 1.256 3.669 1.298 ;
        RECT 3.931 1.256 3.973 1.298 ;
        RECT 1.803 1.282 1.845 1.324 ;
        RECT 1.955 1.282 1.997 1.324 ;
        RECT 0.739 1.292 0.781 1.334 ;
        RECT 3.323 1.3 3.365 1.342 ;
        RECT 0.891 1.306 0.933 1.348 ;
        RECT 2.715 1.312 2.757 1.354 ;
        RECT 3.171 1.312 3.213 1.354 ;
        RECT 3.627 1.348 3.669 1.39 ;
        RECT 3.931 1.348 3.973 1.39 ;
        RECT 3.323 1.392 3.365 1.434 ;
        RECT 0.891 1.398 0.933 1.44 ;
        RECT 3.627 1.44 3.669 1.482 ;
        RECT 3.323 1.484 3.365 1.526 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
        RECT 3.095 1.651 3.137 1.693 ;
        RECT 3.247 1.651 3.289 1.693 ;
        RECT 3.399 1.651 3.441 1.693 ;
        RECT 3.551 1.651 3.593 1.693 ;
        RECT 3.703 1.651 3.745 1.693 ;
        RECT 3.855 1.651 3.897 1.693 ;
        RECT 4.007 1.651 4.049 1.693 ;
        RECT 4.159 1.651 4.201 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 4.256 1.702 ;
        RECT 2.639 1.358 2.689 1.642 ;
        RECT 3.207 1.358 3.257 1.642 ;
        RECT 0.887 1.354 0.937 1.642 ;
        RECT 1.975 1.328 2.025 1.642 ;
        RECT 2.639 1.308 2.777 1.358 ;
        RECT 3.149 1.308 3.257 1.358 ;
        RECT 0.279 1.033 0.329 1.642 ;
        RECT 3.319 0.912 3.369 1.642 ;
        RECT 3.623 0.96 3.673 1.642 ;
        RECT 3.927 1.052 3.977 1.642 ;
        RECT 0.735 1.304 0.937 1.354 ;
        RECT 1.782 1.278 2.025 1.328 ;
        RECT 0.735 1.088 0.785 1.304 ;
        RECT 0.887 1.101 0.937 1.304 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 3.399 -0.021 3.441 0.021 ;
        RECT 3.551 -0.021 3.593 0.021 ;
        RECT 3.703 -0.021 3.745 0.021 ;
        RECT 3.855 -0.021 3.897 0.021 ;
        RECT 4.007 -0.021 4.049 0.021 ;
        RECT 4.159 -0.021 4.201 0.021 ;
        RECT 3.323 0.158 3.365 0.2 ;
        RECT 3.627 0.158 3.669 0.2 ;
        RECT 3.931 0.158 3.973 0.2 ;
        RECT 0.739 0.2 0.781 0.242 ;
        RECT 1.955 0.203 1.997 0.245 ;
        RECT 1.803 0.219 1.845 0.261 ;
        RECT 3.323 0.25 3.365 0.292 ;
        RECT 3.627 0.25 3.669 0.292 ;
        RECT 0.891 0.275 0.933 0.317 ;
        RECT 1.803 0.311 1.845 0.353 ;
        RECT 2.715 0.334 2.757 0.376 ;
        RECT 3.171 0.334 3.213 0.376 ;
        RECT 3.323 0.342 3.365 0.384 ;
        RECT 0.283 0.344 0.325 0.386 ;
        RECT 0.739 0.388 0.781 0.43 ;
        RECT 0.891 0.388 0.933 0.43 ;
      LAYER M1 ;
        RECT 2.695 0.33 3.233 0.38 ;
        RECT 1.799 0.249 1.849 0.373 ;
        RECT 0.735 0.246 0.785 0.45 ;
        RECT 0.887 0.246 0.937 0.45 ;
        RECT 1.799 0.199 2.024 0.249 ;
        RECT 0.586 0.196 0.937 0.246 ;
        RECT 0.279 0.03 0.329 0.419 ;
        RECT 3.319 0.03 3.369 0.408 ;
        RECT 3.167 0.03 3.217 0.33 ;
        RECT 3.623 0.03 3.673 0.319 ;
        RECT 3.927 0.03 3.977 0.22 ;
        RECT 1.799 0.03 1.849 0.199 ;
        RECT 0.586 0.03 0.636 0.196 ;
        RECT 0 -0.03 4.256 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.191 0.299 1.281 0.381 ;
      RECT 0.431 0.988 1.265 1.038 ;
      RECT 1.191 1.038 1.241 1.314 ;
      RECT 1.215 0.381 1.265 0.988 ;
      RECT 0.431 0.779 0.521 0.829 ;
      RECT 0.431 0.579 0.521 0.629 ;
      RECT 0.431 1.038 0.481 1.216 ;
      RECT 0.431 0.829 0.481 0.988 ;
      RECT 0.431 0.455 0.481 0.579 ;
      RECT 0.471 0.629 0.521 0.779 ;
      RECT 2.115 0.23 2.837 0.28 ;
      RECT 2.787 0.088 2.837 0.23 ;
      RECT 1.964 0.314 2.165 0.364 ;
      RECT 1.707 0.54 2.014 0.59 ;
      RECT 2.315 0.178 2.397 0.23 ;
      RECT 2.115 0.28 2.165 0.314 ;
      RECT 1.964 0.364 2.014 0.54 ;
      RECT 1.343 0.64 2.093 0.69 ;
      RECT 1.343 0.434 1.561 0.484 ;
      RECT 1.343 1.158 1.561 1.208 ;
      RECT 1.343 0.355 1.393 0.434 ;
      RECT 1.343 1.208 1.393 1.314 ;
      RECT 1.343 0.69 1.393 1.158 ;
      RECT 1.343 0.484 1.393 0.64 ;
      RECT 3.68 0.604 3.917 0.654 ;
      RECT 2.71 0.494 3.73 0.544 ;
      RECT 3.68 0.544 3.73 0.604 ;
      RECT 3.68 0.654 3.73 0.704 ;
      RECT 3.207 0.704 3.73 0.754 ;
      RECT 2.407 0.438 2.76 0.488 ;
      RECT 2.619 0.699 2.76 0.749 ;
      RECT 2.847 1.208 3.257 1.258 ;
      RECT 2.407 0.488 2.457 1.165 ;
      RECT 3.207 0.754 3.257 1.208 ;
      RECT 2.71 0.544 2.76 0.699 ;
      RECT 2.71 0.488 2.76 0.494 ;
      RECT 1.707 0.758 2.229 0.808 ;
      RECT 2.179 0.587 2.229 0.758 ;
      RECT 1.55 1.001 2.345 1.051 ;
      RECT 2.255 0.371 2.305 0.42 ;
      RECT 2.072 0.42 2.345 0.47 ;
      RECT 2.103 1.166 2.153 1.308 ;
      RECT 2.103 1.308 2.305 1.358 ;
      RECT 2.295 0.47 2.345 1.001 ;
      RECT 2.255 1.051 2.305 1.308 ;
      RECT 2.77 1.521 3.157 1.571 ;
      RECT 1.419 1.478 1.789 1.528 ;
      RECT 1.419 1.528 1.469 1.565 ;
      RECT 1.099 1.526 1.317 1.576 ;
      RECT 1.875 1.428 1.925 1.584 ;
      RECT 1.267 1.428 1.317 1.526 ;
      RECT 1.267 1.378 1.925 1.428 ;
      RECT 0.583 0.618 1.029 0.668 ;
      RECT 0.583 0.668 0.633 0.914 ;
      RECT 0.583 0.422 0.633 0.618 ;
      RECT 1.039 0.518 1.165 0.568 ;
      RECT 1.039 0.768 1.089 0.914 ;
      RECT 1.039 0.718 1.165 0.768 ;
      RECT 1.039 0.394 1.089 0.518 ;
      RECT 1.115 0.568 1.165 0.718 ;
      RECT 2.824 0.604 3.613 0.654 ;
      RECT 2.519 0.588 2.569 0.978 ;
      RECT 2.519 0.538 2.625 0.588 ;
      RECT 2.542 1.027 2.874 1.028 ;
      RECT 2.824 1.028 2.874 1.029 ;
      RECT 2.824 0.654 2.874 0.978 ;
      RECT 2.519 0.978 2.874 1.027 ;
      RECT 2.934 0.709 3.157 0.759 ;
      RECT 2.355 1.272 2.581 1.322 ;
      RECT 2.163 1.522 2.405 1.572 ;
      RECT 2.355 1.322 2.405 1.522 ;
      RECT 2.531 1.149 2.581 1.272 ;
      RECT 2.934 0.759 2.984 1.099 ;
      RECT 2.531 1.099 2.984 1.149 ;
      RECT 0.795 0.096 1.491 0.146 ;
    LAYER CO ;
      RECT 1.195 0.319 1.237 0.361 ;
      RECT 1.347 0.375 1.389 0.417 ;
      RECT 1.727 0.762 1.769 0.804 ;
      RECT 1.879 1.522 1.921 1.564 ;
      RECT 1.195 1.252 1.237 1.294 ;
      RECT 1.043 0.506 1.085 0.548 ;
      RECT 0.435 1.062 0.477 1.104 ;
      RECT 1.043 0.414 1.085 0.456 ;
      RECT 2.107 1.199 2.149 1.241 ;
      RECT 2.107 1.291 2.149 1.333 ;
      RECT 2.867 1.212 2.909 1.254 ;
      RECT 3.703 0.608 3.745 0.65 ;
      RECT 3.855 0.608 3.897 0.65 ;
      RECT 3.399 0.608 3.441 0.65 ;
      RECT 1.043 0.852 1.085 0.894 ;
      RECT 2.259 0.391 2.301 0.433 ;
      RECT 1.347 0.375 1.389 0.417 ;
      RECT 1.195 0.319 1.237 0.361 ;
      RECT 1.195 0.319 1.237 0.361 ;
      RECT 0.587 0.852 0.629 0.894 ;
      RECT 3.095 0.713 3.137 0.755 ;
      RECT 0.435 1.154 0.477 1.196 ;
      RECT 0.435 1.062 0.477 1.104 ;
      RECT 1.499 1.162 1.541 1.204 ;
      RECT 1.347 1.16 1.389 1.202 ;
      RECT 1.119 1.53 1.161 1.572 ;
      RECT 1.727 1.482 1.769 1.524 ;
      RECT 0.587 0.76 0.629 0.802 ;
      RECT 2.031 0.644 2.073 0.686 ;
      RECT 2.259 1.107 2.301 1.149 ;
      RECT 3.095 1.525 3.137 1.567 ;
      RECT 2.183 1.526 2.225 1.568 ;
      RECT 1.271 1.49 1.313 1.532 ;
      RECT 2.791 1.525 2.833 1.567 ;
      RECT 2.639 0.703 2.681 0.745 ;
      RECT 2.867 0.498 2.909 0.54 ;
      RECT 2.411 0.49 2.453 0.532 ;
      RECT 2.183 0.644 2.225 0.686 ;
      RECT 2.791 0.128 2.833 0.17 ;
      RECT 2.335 0.18 2.377 0.222 ;
      RECT 1.727 0.544 1.769 0.586 ;
      RECT 1.499 0.438 1.541 0.48 ;
      RECT 1.423 0.1 1.465 0.142 ;
      RECT 2.943 0.608 2.985 0.65 ;
      RECT 1.575 1.005 1.617 1.047 ;
      RECT 3.551 0.608 3.593 0.65 ;
      RECT 0.815 0.1 0.857 0.142 ;
      RECT 1.119 0.649 1.161 0.691 ;
      RECT 0.435 0.492 0.477 0.534 ;
      RECT 1.195 1.16 1.237 1.202 ;
      RECT 2.335 1.526 2.377 1.568 ;
      RECT 2.563 0.982 2.605 1.024 ;
      RECT 1.043 0.76 1.085 0.802 ;
      RECT 0.815 0.622 0.857 0.664 ;
      RECT 2.259 1.291 2.301 1.333 ;
      RECT 0.435 1.154 0.477 1.196 ;
      RECT 2.411 1.103 2.453 1.145 ;
      RECT 2.107 0.424 2.149 0.466 ;
      RECT 0.967 0.622 1.009 0.664 ;
      RECT 1.347 1.252 1.389 1.294 ;
      RECT 2.563 0.542 2.605 0.584 ;
      RECT 1.879 0.544 1.921 0.586 ;
      RECT 1.423 1.503 1.465 1.545 ;
      RECT 2.259 1.199 2.301 1.241 ;
      RECT 0.587 0.442 0.629 0.484 ;
      RECT 0.587 0.442 0.629 0.484 ;
      RECT 1.271 0.1 1.313 0.142 ;
      RECT 0.587 0.442 0.629 0.484 ;
      RECT 1.347 0.375 1.389 0.417 ;
    LAYER PO ;
      RECT 3.101 1.012 3.131 1.606 ;
      RECT 2.341 0.068 2.371 0.622 ;
      RECT 0.061 0.066 0.091 1.606 ;
      RECT 0.365 0.068 0.395 1.606 ;
      RECT 0.213 0.066 0.243 1.606 ;
      RECT 1.733 0.73 1.763 1.606 ;
      RECT 1.125 0.068 1.155 1.606 ;
      RECT 3.253 0.068 3.283 1.606 ;
      RECT 2.949 0.068 2.979 1.606 ;
      RECT 1.885 0.068 1.915 1.606 ;
      RECT 0.669 0.068 0.699 1.606 ;
      RECT 2.037 0.068 2.067 1.606 ;
      RECT 1.581 0.068 1.611 1.606 ;
      RECT 0.821 0.068 0.851 1.606 ;
      RECT 2.493 0.068 2.523 1.606 ;
      RECT 2.189 0.068 2.219 1.606 ;
      RECT 2.797 0.068 2.827 1.606 ;
      RECT 1.429 0.068 1.459 1.606 ;
      RECT 2.645 0.068 2.675 1.606 ;
      RECT 0.973 0.068 1.003 1.606 ;
      RECT 0.517 0.068 0.547 1.606 ;
      RECT 3.709 0.068 3.739 1.606 ;
      RECT 3.405 0.068 3.435 1.606 ;
      RECT 1.277 0.068 1.307 0.542 ;
      RECT 1.277 0.99 1.307 1.606 ;
      RECT 3.101 0.068 3.131 0.787 ;
      RECT 4.165 0.068 4.195 1.606 ;
      RECT 1.733 0.068 1.763 0.618 ;
      RECT 3.557 0.068 3.587 1.606 ;
      RECT 2.341 0.882 2.371 1.606 ;
      RECT 4.013 0.068 4.043 1.606 ;
      RECT 3.861 0.068 3.891 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 4.371 1.773 ;
  END
END DFFX2_RVT

MACRO DFFARX2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 4.56 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.684 0.401 0.726 ;
      LAYER M1 ;
        RECT 0.249 0.68 0.421 0.73 ;
        RECT 0.249 0.553 0.359 0.68 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 ;
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 1.53 0.705 1.572 ;
      LAYER M1 ;
        RECT 0.553 1.424 0.725 1.576 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 2.791 0.118 2.833 0.16 ;
        RECT 1.727 0.122 1.769 0.164 ;
      LAYER M1 ;
        RECT 1.723 0.138 1.879 0.207 ;
        RECT 2.771 0.138 2.853 0.174 ;
        RECT 1.723 0.088 2.853 0.138 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0441 ;
  END RSTB
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.779 0.195 3.821 0.237 ;
        RECT 3.779 0.287 3.821 0.329 ;
        RECT 3.779 0.932 3.821 0.974 ;
        RECT 3.779 1.024 3.821 1.066 ;
        RECT 3.779 1.116 3.821 1.158 ;
        RECT 3.779 1.208 3.821 1.25 ;
        RECT 3.779 1.3 3.821 1.342 ;
        RECT 3.779 1.392 3.821 1.434 ;
        RECT 3.779 1.484 3.821 1.526 ;
      LAYER M1 ;
        RECT 3.775 0.854 3.825 1.546 ;
        RECT 3.775 0.804 4.321 0.854 ;
        RECT 4.271 0.511 4.321 0.804 ;
        RECT 4.201 0.444 4.321 0.511 ;
        RECT 3.775 0.394 4.321 0.444 ;
        RECT 3.775 0.148 3.825 0.394 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 4.083 0.195 4.125 0.237 ;
        RECT 4.083 1.024 4.125 1.066 ;
        RECT 4.083 1.116 4.125 1.158 ;
        RECT 4.083 1.208 4.125 1.25 ;
        RECT 4.083 1.3 4.125 1.342 ;
        RECT 4.083 1.392 4.125 1.434 ;
        RECT 4.083 1.484 4.125 1.526 ;
      LAYER M1 ;
        RECT 4.079 0.968 4.129 1.546 ;
        RECT 4.079 0.918 4.445 0.968 ;
        RECT 4.395 0.32 4.445 0.918 ;
        RECT 4.079 0.27 4.445 0.32 ;
        RECT 4.079 0.148 4.129 0.27 ;
        RECT 4.395 0.207 4.445 0.27 ;
        RECT 4.353 0.097 4.463 0.207 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 3.627 0.932 3.669 0.974 ;
        RECT 3.931 0.98 3.973 1.022 ;
        RECT 3.627 1.024 3.669 1.066 ;
        RECT 0.283 1.062 0.325 1.104 ;
        RECT 3.931 1.072 3.973 1.114 ;
        RECT 4.235 1.072 4.277 1.114 ;
        RECT 3.627 1.116 3.669 1.158 ;
        RECT 0.739 1.118 0.781 1.16 ;
        RECT 0.891 1.132 0.933 1.174 ;
        RECT 0.283 1.154 0.325 1.196 ;
        RECT 3.931 1.164 3.973 1.206 ;
        RECT 4.235 1.164 4.277 1.206 ;
        RECT 3.627 1.208 3.669 1.25 ;
        RECT 0.739 1.21 0.781 1.252 ;
        RECT 0.891 1.224 0.933 1.266 ;
        RECT 3.931 1.256 3.973 1.298 ;
        RECT 4.235 1.256 4.277 1.298 ;
        RECT 1.955 1.282 1.997 1.324 ;
        RECT 2.107 1.282 2.149 1.324 ;
        RECT 3.627 1.3 3.669 1.342 ;
        RECT 0.739 1.302 0.781 1.344 ;
        RECT 2.867 1.312 2.909 1.354 ;
        RECT 3.475 1.312 3.517 1.354 ;
        RECT 0.891 1.316 0.933 1.358 ;
        RECT 3.931 1.348 3.973 1.39 ;
        RECT 4.235 1.348 4.277 1.39 ;
        RECT 3.627 1.392 3.669 1.434 ;
        RECT 3.931 1.44 3.973 1.482 ;
        RECT 3.627 1.484 3.669 1.526 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
        RECT 3.095 1.651 3.137 1.693 ;
        RECT 3.247 1.651 3.289 1.693 ;
        RECT 3.399 1.651 3.441 1.693 ;
        RECT 3.551 1.651 3.593 1.693 ;
        RECT 3.703 1.651 3.745 1.693 ;
        RECT 3.855 1.651 3.897 1.693 ;
        RECT 4.007 1.651 4.049 1.693 ;
        RECT 4.159 1.651 4.201 1.693 ;
        RECT 4.311 1.651 4.353 1.693 ;
        RECT 4.463 1.651 4.505 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 4.56 1.702 ;
        RECT 0.887 1.364 0.937 1.642 ;
        RECT 3.511 1.358 3.561 1.642 ;
        RECT 2.127 1.328 2.177 1.642 ;
        RECT 0.279 1.033 0.329 1.642 ;
        RECT 3.623 0.912 3.673 1.642 ;
        RECT 3.927 0.96 3.977 1.642 ;
        RECT 4.231 1.052 4.281 1.642 ;
        RECT 0.735 1.314 0.937 1.364 ;
        RECT 2.834 1.308 3.561 1.358 ;
        RECT 1.934 1.278 2.177 1.328 ;
        RECT 0.735 1.098 0.785 1.314 ;
        RECT 0.887 1.111 0.937 1.314 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 3.399 -0.021 3.441 0.021 ;
        RECT 3.551 -0.021 3.593 0.021 ;
        RECT 3.703 -0.021 3.745 0.021 ;
        RECT 3.855 -0.021 3.897 0.021 ;
        RECT 4.007 -0.021 4.049 0.021 ;
        RECT 4.159 -0.021 4.201 0.021 ;
        RECT 4.311 -0.021 4.353 0.021 ;
        RECT 4.463 -0.021 4.505 0.021 ;
        RECT 3.627 0.158 3.669 0.2 ;
        RECT 3.931 0.158 3.973 0.2 ;
        RECT 4.235 0.158 4.277 0.2 ;
        RECT 0.739 0.2 0.781 0.242 ;
        RECT 2.107 0.203 2.149 0.245 ;
        RECT 3.627 0.25 3.669 0.292 ;
        RECT 3.931 0.25 3.973 0.292 ;
        RECT 0.891 0.275 0.933 0.317 ;
        RECT 1.955 0.307 1.997 0.349 ;
        RECT 3.019 0.334 3.061 0.376 ;
        RECT 3.475 0.334 3.517 0.376 ;
        RECT 3.627 0.342 3.669 0.384 ;
        RECT 0.283 0.344 0.325 0.386 ;
        RECT 0.739 0.388 0.781 0.43 ;
        RECT 0.891 0.388 0.933 0.43 ;
        RECT 1.955 0.399 1.997 0.441 ;
      LAYER M1 ;
        RECT 1.951 0.337 2.001 0.461 ;
        RECT 2.999 0.33 3.537 0.38 ;
        RECT 1.541 0.287 2.001 0.337 ;
        RECT 1.951 0.249 2.001 0.287 ;
        RECT 0.735 0.246 0.785 0.45 ;
        RECT 0.887 0.246 0.937 0.45 ;
        RECT 1.951 0.199 2.176 0.249 ;
        RECT 0.586 0.196 0.937 0.246 ;
        RECT 0.279 0.03 0.329 0.419 ;
        RECT 3.623 0.03 3.673 0.408 ;
        RECT 3.471 0.03 3.521 0.33 ;
        RECT 3.927 0.03 3.977 0.319 ;
        RECT 1.541 0.03 1.591 0.287 ;
        RECT 4.231 0.03 4.281 0.22 ;
        RECT 0.586 0.03 0.636 0.196 ;
        RECT 0 -0.03 4.56 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 2.715 0.982 2.757 1.024 ;
      RECT 1.043 0.76 1.085 0.802 ;
      RECT 2.563 1.103 2.605 1.145 ;
      RECT 3.171 1.212 3.213 1.254 ;
      RECT 0.967 0.622 1.009 0.664 ;
      RECT 1.195 0.319 1.237 0.361 ;
      RECT 1.347 0.375 1.389 0.417 ;
      RECT 1.879 0.79 1.921 0.832 ;
      RECT 3.171 0.508 3.213 0.55 ;
      RECT 3.019 0.982 3.061 1.024 ;
      RECT 2.031 1.522 2.073 1.564 ;
      RECT 1.195 1.252 1.237 1.294 ;
      RECT 1.043 0.506 1.085 0.548 ;
      RECT 0.435 1.062 0.477 1.104 ;
      RECT 1.043 0.414 1.085 0.456 ;
      RECT 3.399 0.713 3.441 0.755 ;
      RECT 3.247 0.608 3.289 0.65 ;
      RECT 1.271 0.1 1.313 0.142 ;
      RECT 1.119 1.53 1.161 1.572 ;
      RECT 1.423 0.1 1.465 0.142 ;
      RECT 2.259 1.164 2.301 1.206 ;
      RECT 1.043 0.852 1.085 0.894 ;
      RECT 2.411 0.391 2.453 0.433 ;
      RECT 3.399 1.432 3.441 1.474 ;
      RECT 3.855 0.608 3.897 0.65 ;
      RECT 3.703 0.608 3.745 0.65 ;
      RECT 0.587 0.442 0.629 0.484 ;
      RECT 0.587 0.442 0.629 0.484 ;
      RECT 0.587 0.442 0.629 0.484 ;
      RECT 1.347 0.375 1.389 0.417 ;
      RECT 1.347 0.375 1.389 0.417 ;
      RECT 1.195 0.319 1.237 0.361 ;
      RECT 1.195 0.319 1.237 0.361 ;
      RECT 0.587 0.852 0.629 0.894 ;
      RECT 4.007 0.608 4.049 0.65 ;
      RECT 0.435 1.154 0.477 1.196 ;
      RECT 0.435 1.062 0.477 1.104 ;
      RECT 3.855 0.608 3.897 0.65 ;
      RECT 1.651 1.162 1.693 1.204 ;
      RECT 1.347 1.16 1.389 1.202 ;
      RECT 0.815 0.1 0.857 0.142 ;
      RECT 1.879 1.482 1.921 1.524 ;
      RECT 4.159 0.608 4.201 0.65 ;
      RECT 0.587 0.76 0.629 0.802 ;
      RECT 2.183 0.644 2.225 0.686 ;
      RECT 2.411 1.107 2.453 1.149 ;
      RECT 2.259 1.282 2.301 1.324 ;
      RECT 3.703 0.608 3.745 0.65 ;
      RECT 2.335 1.532 2.377 1.574 ;
      RECT 1.271 1.49 1.313 1.532 ;
      RECT 3.095 1.433 3.137 1.475 ;
      RECT 1.499 1.282 1.541 1.324 ;
      RECT 2.943 0.77 2.985 0.812 ;
      RECT 2.563 0.49 2.605 0.532 ;
      RECT 3.095 0.12 3.137 0.162 ;
      RECT 2.487 0.19 2.529 0.232 ;
      RECT 1.879 0.544 1.921 0.586 ;
      RECT 1.499 0.438 1.541 0.48 ;
      RECT 2.335 0.641 2.377 0.683 ;
      RECT 1.575 1.005 1.617 1.047 ;
      RECT 1.803 1.282 1.845 1.324 ;
      RECT 1.119 0.649 1.161 0.691 ;
      RECT 0.435 0.492 0.477 0.534 ;
      RECT 1.195 1.16 1.237 1.202 ;
      RECT 2.487 1.532 2.529 1.574 ;
      RECT 0.815 0.622 0.857 0.664 ;
      RECT 2.411 1.291 2.453 1.333 ;
      RECT 0.435 1.154 0.477 1.196 ;
      RECT 2.259 0.424 2.301 0.466 ;
      RECT 1.347 1.252 1.389 1.294 ;
      RECT 2.715 0.542 2.757 0.584 ;
      RECT 2.031 0.544 2.073 0.586 ;
      RECT 1.423 1.503 1.465 1.545 ;
      RECT 2.411 1.199 2.453 1.241 ;
    LAYER M1 ;
      RECT 1.191 0.299 1.281 0.381 ;
      RECT 1.191 1.038 1.241 1.314 ;
      RECT 0.431 0.988 1.265 1.038 ;
      RECT 1.215 0.381 1.265 0.988 ;
      RECT 0.431 0.779 0.521 0.829 ;
      RECT 0.431 0.579 0.521 0.629 ;
      RECT 0.431 1.038 0.481 1.216 ;
      RECT 0.431 0.829 0.481 0.988 ;
      RECT 0.431 0.455 0.481 0.579 ;
      RECT 0.471 0.629 0.521 0.779 ;
      RECT 2.249 0.23 3.141 0.28 ;
      RECT 3.091 0.088 3.141 0.23 ;
      RECT 2.098 0.314 2.299 0.364 ;
      RECT 1.859 0.54 2.148 0.59 ;
      RECT 2.467 0.188 2.549 0.23 ;
      RECT 2.249 0.28 2.299 0.314 ;
      RECT 2.098 0.364 2.148 0.54 ;
      RECT 1.343 0.64 2.245 0.69 ;
      RECT 1.343 0.434 1.561 0.484 ;
      RECT 1.343 1.158 1.713 1.208 ;
      RECT 1.343 0.355 1.393 0.434 ;
      RECT 1.343 1.208 1.393 1.314 ;
      RECT 1.343 0.69 1.393 1.158 ;
      RECT 1.343 0.484 1.393 0.64 ;
      RECT 3.984 0.604 4.221 0.654 ;
      RECT 2.862 0.504 4.034 0.554 ;
      RECT 3.984 0.503 4.034 0.504 ;
      RECT 3.984 0.554 4.034 0.604 ;
      RECT 3.984 0.654 4.034 0.704 ;
      RECT 3.511 0.704 4.034 0.754 ;
      RECT 2.559 0.438 2.912 0.488 ;
      RECT 3.151 1.208 3.561 1.258 ;
      RECT 2.559 0.488 2.609 1.165 ;
      RECT 2.862 0.766 3.005 0.816 ;
      RECT 3.511 0.754 3.561 1.208 ;
      RECT 2.862 0.554 2.912 0.766 ;
      RECT 2.862 0.488 2.912 0.504 ;
      RECT 1.859 0.786 2.381 0.836 ;
      RECT 2.331 0.621 2.381 0.786 ;
      RECT 2.407 0.509 2.497 0.559 ;
      RECT 1.55 1.001 2.497 1.051 ;
      RECT 2.224 0.42 2.457 0.47 ;
      RECT 2.255 1.308 2.457 1.358 ;
      RECT 2.447 0.559 2.497 1.001 ;
      RECT 2.407 0.47 2.457 0.509 ;
      RECT 2.407 0.371 2.457 0.42 ;
      RECT 2.255 1.101 2.305 1.308 ;
      RECT 2.407 1.051 2.457 1.308 ;
      RECT 0.781 0.096 1.491 0.146 ;
      RECT 3.055 0.604 3.917 0.654 ;
      RECT 2.694 0.978 3.105 1.028 ;
      RECT 2.694 0.538 2.801 0.588 ;
      RECT 3.055 0.654 3.105 0.978 ;
      RECT 2.694 0.588 2.744 0.978 ;
      RECT 1.419 1.478 1.941 1.528 ;
      RECT 1.419 1.528 1.469 1.565 ;
      RECT 1.087 1.526 1.317 1.576 ;
      RECT 2.027 1.428 2.077 1.584 ;
      RECT 1.267 1.428 1.317 1.526 ;
      RECT 1.267 1.378 2.077 1.428 ;
      RECT 0.583 0.618 1.029 0.668 ;
      RECT 0.583 0.668 0.633 0.914 ;
      RECT 0.583 0.422 0.633 0.618 ;
      RECT 1.039 0.518 1.165 0.568 ;
      RECT 1.039 0.768 1.089 0.914 ;
      RECT 1.039 0.718 1.165 0.768 ;
      RECT 1.039 0.394 1.089 0.518 ;
      RECT 1.115 0.568 1.165 0.718 ;
      RECT 3.074 1.429 3.461 1.479 ;
      RECT 3.238 0.709 3.461 0.759 ;
      RECT 3.238 0.759 3.288 1.099 ;
      RECT 2.683 1.099 3.288 1.149 ;
      RECT 2.507 1.272 2.733 1.322 ;
      RECT 2.315 1.528 2.557 1.578 ;
      RECT 2.507 1.322 2.557 1.528 ;
      RECT 2.683 1.149 2.733 1.272 ;
      RECT 1.479 1.278 1.865 1.328 ;
    LAYER PO ;
      RECT 2.493 0.068 2.523 0.632 ;
      RECT 3.253 0.068 3.283 1.606 ;
      RECT 0.061 0.066 0.091 1.606 ;
      RECT 0.365 0.068 0.395 1.606 ;
      RECT 0.213 0.066 0.243 1.606 ;
      RECT 1.885 0.758 1.915 1.606 ;
      RECT 1.125 0.068 1.155 1.606 ;
      RECT 3.557 0.068 3.587 1.606 ;
      RECT 2.949 0.068 2.979 1.606 ;
      RECT 2.037 0.068 2.067 1.606 ;
      RECT 0.669 0.068 0.699 1.606 ;
      RECT 1.733 0.068 1.763 1.606 ;
      RECT 0.821 0.068 0.851 1.606 ;
      RECT 2.645 0.068 2.675 1.606 ;
      RECT 2.341 0.068 2.371 1.606 ;
      RECT 3.101 0.068 3.131 1.606 ;
      RECT 1.429 0.068 1.459 1.606 ;
      RECT 2.797 0.068 2.827 1.606 ;
      RECT 0.973 0.068 1.003 1.606 ;
      RECT 1.581 0.068 1.611 1.606 ;
      RECT 0.517 0.068 0.547 1.606 ;
      RECT 1.277 0.068 1.307 0.542 ;
      RECT 1.277 0.99 1.307 1.606 ;
      RECT 3.405 1.012 3.435 1.606 ;
      RECT 3.709 0.068 3.739 1.606 ;
      RECT 2.189 0.068 2.219 1.606 ;
      RECT 3.861 0.068 3.891 1.606 ;
      RECT 4.013 0.068 4.043 1.606 ;
      RECT 4.469 0.068 4.499 1.606 ;
      RECT 1.885 0.068 1.915 0.618 ;
      RECT 3.405 0.068 3.435 0.787 ;
      RECT 2.493 0.882 2.523 1.606 ;
      RECT 4.165 0.068 4.195 1.606 ;
      RECT 4.317 0.068 4.347 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 4.675 1.773 ;
  END
END DFFARX2_RVT

MACRO DFFSSRX2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 4.56 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.881 0.857 0.923 ;
      LAYER M1 ;
        RECT 0.795 0.857 0.967 0.977 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 ;
  END D
  PIN SETB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.207 0.705 0.249 0.747 ;
      LAYER M1 ;
        RECT 0.097 0.751 0.207 0.825 ;
        RECT 0.097 0.701 0.269 0.751 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 ;
  END SETB
  PIN RSTB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.205 0.401 0.247 ;
        RECT 0.511 0.205 0.553 0.247 ;
      LAYER M1 ;
        RECT 0.249 0.201 0.573 0.251 ;
        RECT 0.249 0.097 0.359 0.201 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 ;
  END RSTB
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.119 1.532 1.161 1.574 ;
      LAYER M1 ;
        RECT 1.009 1.465 1.181 1.576 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 4.083 0.195 4.125 0.237 ;
        RECT 4.083 1.024 4.125 1.066 ;
        RECT 4.083 1.116 4.125 1.158 ;
        RECT 4.083 1.208 4.125 1.25 ;
        RECT 4.083 1.3 4.125 1.342 ;
        RECT 4.083 1.392 4.125 1.434 ;
        RECT 4.083 1.484 4.125 1.526 ;
      LAYER M1 ;
        RECT 4.079 0.968 4.129 1.546 ;
        RECT 4.079 0.918 4.445 0.968 ;
        RECT 4.395 0.359 4.445 0.918 ;
        RECT 4.353 0.32 4.463 0.359 ;
        RECT 4.079 0.27 4.463 0.32 ;
        RECT 4.079 0.148 4.129 0.27 ;
        RECT 4.353 0.217 4.463 0.27 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.779 0.195 3.821 0.237 ;
        RECT 3.779 0.287 3.821 0.329 ;
        RECT 3.779 0.932 3.821 0.974 ;
        RECT 3.779 1.024 3.821 1.066 ;
        RECT 3.779 1.116 3.821 1.158 ;
        RECT 3.779 1.208 3.821 1.25 ;
        RECT 3.779 1.3 3.821 1.342 ;
        RECT 3.779 1.392 3.821 1.434 ;
        RECT 3.779 1.484 3.821 1.526 ;
      LAYER M1 ;
        RECT 3.775 0.854 3.825 1.546 ;
        RECT 3.775 0.804 4.321 0.854 ;
        RECT 4.271 0.511 4.321 0.804 ;
        RECT 4.201 0.444 4.321 0.511 ;
        RECT 3.775 0.401 4.321 0.444 ;
        RECT 3.775 0.394 4.283 0.401 ;
        RECT 3.775 0.148 3.825 0.394 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 3.627 0.932 3.669 0.974 ;
        RECT 0.131 0.95 0.173 0.992 ;
        RECT 3.931 0.98 3.973 1.022 ;
        RECT 0.435 1 0.477 1.042 ;
        RECT 3.627 1.024 3.669 1.066 ;
        RECT 0.131 1.042 0.173 1.084 ;
        RECT 3.931 1.072 3.973 1.114 ;
        RECT 4.235 1.072 4.277 1.114 ;
        RECT 0.435 1.092 0.477 1.134 ;
        RECT 3.627 1.116 3.669 1.158 ;
        RECT 2.107 1.12 2.149 1.162 ;
        RECT 0.131 1.134 0.173 1.176 ;
        RECT 3.931 1.164 3.973 1.206 ;
        RECT 4.235 1.164 4.277 1.206 ;
        RECT 0.435 1.184 0.477 1.226 ;
        RECT 3.627 1.208 3.669 1.25 ;
        RECT 2.107 1.212 2.149 1.254 ;
        RECT 0.131 1.226 0.173 1.268 ;
        RECT 3.475 1.236 3.517 1.278 ;
        RECT 3.931 1.256 3.973 1.298 ;
        RECT 4.235 1.256 4.277 1.298 ;
        RECT 0.435 1.276 0.477 1.318 ;
        RECT 3.627 1.3 3.669 1.342 ;
        RECT 2.107 1.304 2.149 1.346 ;
        RECT 0.131 1.318 0.173 1.36 ;
        RECT 1.195 1.32 1.237 1.362 ;
        RECT 3.475 1.328 3.517 1.37 ;
        RECT 2.259 1.336 2.301 1.378 ;
        RECT 3.931 1.348 3.973 1.39 ;
        RECT 4.235 1.348 4.277 1.39 ;
        RECT 3.627 1.392 3.669 1.434 ;
        RECT 3.019 1.42 3.061 1.462 ;
        RECT 3.475 1.42 3.517 1.462 ;
        RECT 2.259 1.428 2.301 1.47 ;
        RECT 3.931 1.44 3.973 1.482 ;
        RECT 3.627 1.484 3.669 1.526 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
        RECT 3.095 1.651 3.137 1.693 ;
        RECT 3.247 1.651 3.289 1.693 ;
        RECT 3.399 1.651 3.441 1.693 ;
        RECT 3.551 1.651 3.593 1.693 ;
        RECT 3.703 1.651 3.745 1.693 ;
        RECT 3.855 1.651 3.897 1.693 ;
        RECT 4.007 1.651 4.049 1.693 ;
        RECT 4.159 1.651 4.201 1.693 ;
        RECT 4.311 1.651 4.353 1.693 ;
        RECT 4.463 1.651 4.505 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 4.56 1.702 ;
        RECT 3.511 1.466 3.561 1.642 ;
        RECT 2.999 1.416 3.561 1.466 ;
        RECT 1.253 1.366 1.303 1.642 ;
        RECT 2.255 1.366 2.305 1.642 ;
        RECT 0.127 1.346 0.177 1.642 ;
        RECT 1.153 1.316 1.303 1.366 ;
        RECT 2.103 1.316 2.305 1.366 ;
        RECT 3.623 0.912 3.673 1.642 ;
        RECT 3.927 0.96 3.977 1.642 ;
        RECT 4.231 1.052 4.281 1.642 ;
        RECT 3.471 1.192 3.521 1.416 ;
        RECT 0.127 1.296 0.481 1.346 ;
        RECT 2.103 1.1 2.153 1.316 ;
        RECT 0.127 0.93 0.177 1.296 ;
        RECT 0.431 0.98 0.481 1.296 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 3.399 -0.021 3.441 0.021 ;
        RECT 3.551 -0.021 3.593 0.021 ;
        RECT 3.703 -0.021 3.745 0.021 ;
        RECT 3.855 -0.021 3.897 0.021 ;
        RECT 4.007 -0.021 4.049 0.021 ;
        RECT 4.159 -0.021 4.201 0.021 ;
        RECT 4.311 -0.021 4.353 0.021 ;
        RECT 4.463 -0.021 4.505 0.021 ;
        RECT 3.627 0.158 3.669 0.2 ;
        RECT 3.931 0.158 3.973 0.2 ;
        RECT 4.235 0.158 4.277 0.2 ;
        RECT 3.019 0.208 3.061 0.25 ;
        RECT 3.475 0.247 3.517 0.289 ;
        RECT 3.627 0.25 3.669 0.292 ;
        RECT 3.931 0.25 3.973 0.292 ;
        RECT 2.107 0.321 2.149 0.363 ;
        RECT 2.259 0.321 2.301 0.363 ;
        RECT 3.475 0.339 3.517 0.381 ;
        RECT 3.627 0.342 3.669 0.384 ;
        RECT 0.131 0.359 0.173 0.401 ;
        RECT 0.435 0.375 0.477 0.417 ;
        RECT 1.195 0.396 1.237 0.438 ;
        RECT 2.107 0.413 2.149 0.455 ;
        RECT 2.259 0.413 2.301 0.455 ;
        RECT 0.131 0.451 0.173 0.493 ;
        RECT 0.435 0.467 0.477 0.509 ;
        RECT 1.195 0.488 1.237 0.53 ;
      LAYER M1 ;
        RECT 0.431 0.405 0.481 0.529 ;
        RECT 0.127 0.405 0.177 0.513 ;
        RECT 0.127 0.355 0.481 0.405 ;
        RECT 1.191 0.351 1.241 0.576 ;
        RECT 2.103 0.351 2.153 0.475 ;
        RECT 2.255 0.351 2.305 0.475 ;
        RECT 1.191 0.301 2.305 0.351 ;
        RECT 2.975 0.204 3.081 0.254 ;
        RECT 3.623 0.03 3.673 0.408 ;
        RECT 3.471 0.03 3.521 0.401 ;
        RECT 0.127 0.03 0.177 0.355 ;
        RECT 3.927 0.03 3.977 0.319 ;
        RECT 1.875 0.03 1.925 0.301 ;
        RECT 4.231 0.03 4.281 0.22 ;
        RECT 2.975 0.03 3.025 0.204 ;
        RECT 0 -0.03 4.56 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 3.703 0.608 3.745 0.65 ;
      RECT 3.703 0.608 3.745 0.65 ;
      RECT 3.855 0.608 3.897 0.65 ;
      RECT 0.283 1.092 0.325 1.134 ;
      RECT 0.283 1 0.325 1.042 ;
      RECT 2.411 1.104 2.453 1.146 ;
      RECT 1.347 0.45 1.389 0.492 ;
      RECT 0.587 0.305 0.629 0.347 ;
      RECT 1.043 0.814 1.085 0.856 ;
      RECT 0.283 1.092 0.325 1.134 ;
      RECT 1.347 0.906 1.389 0.948 ;
      RECT 2.867 0.308 2.909 0.35 ;
      RECT 0.587 1.184 0.629 1.226 ;
      RECT 1.499 0.45 1.541 0.492 ;
      RECT 2.563 1.213 2.605 1.255 ;
      RECT 1.727 1.421 1.769 1.463 ;
      RECT 1.651 1.082 1.693 1.124 ;
      RECT 0.587 1.092 0.629 1.134 ;
      RECT 1.043 0.998 1.085 1.04 ;
      RECT 2.639 1.532 2.681 1.574 ;
      RECT 1.499 1.082 1.541 1.124 ;
      RECT 2.715 1.199 2.757 1.241 ;
      RECT 0.511 0.848 0.553 0.89 ;
      RECT 1.499 0.45 1.541 0.492 ;
      RECT 2.563 0.32 2.605 0.362 ;
      RECT 1.651 0.45 1.693 0.492 ;
      RECT 3.855 0.608 3.897 0.65 ;
      RECT 4.007 0.608 4.049 0.65 ;
      RECT 4.159 0.608 4.201 0.65 ;
      RECT 2.639 0.155 2.681 0.197 ;
      RECT 3.171 1.22 3.213 1.262 ;
      RECT 2.791 0.108 2.833 0.15 ;
      RECT 1.043 1.09 1.085 1.132 ;
      RECT 0.739 1.092 0.781 1.134 ;
      RECT 1.347 0.45 1.389 0.492 ;
      RECT 2.031 0.155 2.073 0.197 ;
      RECT 1.347 0.906 1.389 0.948 ;
      RECT 1.423 1.532 1.465 1.574 ;
      RECT 2.715 0.412 2.757 0.454 ;
      RECT 0.663 1.453 0.705 1.495 ;
      RECT 2.715 0.32 2.757 0.362 ;
      RECT 1.043 0.998 1.085 1.04 ;
      RECT 0.891 0.305 0.933 0.347 ;
      RECT 0.587 1.092 0.629 1.134 ;
      RECT 1.347 0.814 1.389 0.856 ;
      RECT 0.587 1.184 0.629 1.226 ;
      RECT 0.739 0.447 0.781 0.489 ;
      RECT 2.563 1.305 2.605 1.347 ;
      RECT 0.663 0.577 0.705 0.619 ;
      RECT 1.803 1.092 1.845 1.134 ;
      RECT 3.171 0.481 3.213 0.523 ;
      RECT 0.739 1.184 0.781 1.226 ;
      RECT 1.651 0.99 1.693 1.032 ;
      RECT 1.651 0.45 1.693 0.492 ;
      RECT 0.967 0.108 1.009 0.15 ;
      RECT 0.739 1.184 0.781 1.226 ;
      RECT 1.347 0.998 1.389 1.04 ;
      RECT 0.891 1.32 0.933 1.362 ;
      RECT 3.247 0.108 3.289 0.15 ;
      RECT 1.043 0.906 1.085 0.948 ;
      RECT 2.563 0.412 2.605 0.454 ;
      RECT 1.499 0.99 1.541 1.032 ;
      RECT 2.943 0.658 2.985 0.7 ;
      RECT 2.031 0.998 2.073 1.04 ;
      RECT 1.423 0.63 1.465 0.672 ;
      RECT 3.399 1.532 3.441 1.574 ;
      RECT 0.739 1.092 0.781 1.134 ;
      RECT 0.587 1.276 0.629 1.318 ;
      RECT 0.283 1.184 0.325 1.226 ;
      RECT 1.347 0.814 1.389 0.856 ;
      RECT 2.031 1.421 2.073 1.463 ;
      RECT 0.283 1.184 0.325 1.226 ;
      RECT 2.335 0.577 2.377 0.619 ;
      RECT 2.563 1.121 2.605 1.163 ;
      RECT 1.651 0.45 1.693 0.492 ;
      RECT 2.487 1.532 2.529 1.574 ;
      RECT 1.575 1.532 1.617 1.574 ;
      RECT 2.791 1.532 2.833 1.574 ;
      RECT 1.043 0.814 1.085 0.856 ;
      RECT 0.283 0.475 0.325 0.517 ;
      RECT 2.411 0.32 2.453 0.362 ;
      RECT 1.347 0.998 1.389 1.04 ;
      RECT 1.803 1.184 1.845 1.226 ;
      RECT 1.651 1.174 1.693 1.216 ;
      RECT 1.043 0.906 1.085 0.948 ;
      RECT 1.575 0.155 1.617 0.197 ;
      RECT 1.043 0.513 1.085 0.555 ;
      RECT 2.411 0.412 2.453 0.454 ;
      RECT 1.347 0.45 1.389 0.492 ;
      RECT 1.043 0.421 1.085 0.463 ;
      RECT 1.499 0.45 1.541 0.492 ;
      RECT 1.879 0.777 1.921 0.819 ;
      RECT 0.587 1 0.629 1.042 ;
      RECT 3.399 0.681 3.441 0.723 ;
      RECT 0.587 1 0.629 1.042 ;
      RECT 0.967 0.63 1.009 0.672 ;
      RECT 1.347 1.09 1.389 1.132 ;
      RECT 3.247 0.581 3.289 0.623 ;
      RECT 1.727 0.108 1.769 0.15 ;
      RECT 1.803 0.45 1.845 0.492 ;
      RECT 1.499 1.174 1.541 1.216 ;
      RECT 2.031 0.677 2.073 0.719 ;
      RECT 2.867 1.104 2.909 1.146 ;
      RECT 1.271 0.63 1.313 0.672 ;
      RECT 0.359 1.453 0.401 1.495 ;
      RECT 3.095 0.108 3.137 0.15 ;
      RECT 0.283 1 0.325 1.042 ;
    LAYER M1 ;
      RECT 1.343 0.726 1.445 0.776 ;
      RECT 1.327 0.446 1.445 0.496 ;
      RECT 1.395 0.626 1.485 0.676 ;
      RECT 1.343 0.776 1.393 1.152 ;
      RECT 1.395 0.676 1.445 0.726 ;
      RECT 1.395 0.496 1.445 0.626 ;
      RECT 3.66 0.604 3.917 0.654 ;
      RECT 3.127 0.477 3.71 0.527 ;
      RECT 3.66 0.527 3.71 0.604 ;
      RECT 2.711 1.216 3.257 1.266 ;
      RECT 2.711 0.3 2.761 1.216 ;
      RECT 2.923 0.654 3.177 0.677 ;
      RECT 3.127 0.704 3.257 0.727 ;
      RECT 2.923 0.677 3.257 0.704 ;
      RECT 3.207 0.727 3.257 1.216 ;
      RECT 3.127 0.527 3.177 0.654 ;
      RECT 1.854 0.773 2.609 0.823 ;
      RECT 2.559 0.3 2.609 0.452 ;
      RECT 2.407 0.3 2.457 0.452 ;
      RECT 2.407 0.452 2.609 0.502 ;
      RECT 2.407 0.823 2.457 1.166 ;
      RECT 2.559 0.823 2.609 1.38 ;
      RECT 2.559 0.502 2.609 0.773 ;
      RECT 0.735 1.202 1.545 1.252 ;
      RECT 1.495 0.726 1.585 0.776 ;
      RECT 1.495 0.526 1.585 0.576 ;
      RECT 1.495 0.776 1.545 1.202 ;
      RECT 1.495 0.43 1.545 0.526 ;
      RECT 1.535 0.576 1.585 0.726 ;
      RECT 0.695 0.752 0.854 0.802 ;
      RECT 0.719 0.443 0.854 0.493 ;
      RECT 0.804 0.493 0.854 0.752 ;
      RECT 0.695 1.047 0.785 1.097 ;
      RECT 0.695 0.802 0.745 1.047 ;
      RECT 0.735 1.097 0.785 1.202 ;
      RECT 2.011 0.154 2.755 0.201 ;
      RECT 2.705 0.104 2.853 0.151 ;
      RECT 2.011 0.151 2.853 0.154 ;
      RECT 2.659 1.316 3.421 1.366 ;
      RECT 3.371 0.677 3.461 0.727 ;
      RECT 3.371 0.727 3.421 1.316 ;
      RECT 2.415 1.528 2.709 1.578 ;
      RECT 2.251 1.216 2.465 1.266 ;
      RECT 2.011 0.994 2.301 1.044 ;
      RECT 2.659 1.366 2.709 1.528 ;
      RECT 2.415 1.266 2.465 1.528 ;
      RECT 2.251 1.044 2.301 1.216 ;
      RECT 1.647 0.573 2.397 0.623 ;
      RECT 1.647 1.196 1.849 1.246 ;
      RECT 1.799 1.072 1.849 1.196 ;
      RECT 1.799 0.43 1.849 0.573 ;
      RECT 1.647 0.623 1.697 1.196 ;
      RECT 1.647 0.43 1.697 0.573 ;
      RECT 0.339 1.449 0.725 1.499 ;
      RECT 3.075 0.104 3.309 0.154 ;
      RECT 2.823 0.304 3.226 0.354 ;
      RECT 3.176 0.154 3.226 0.304 ;
      RECT 2.823 0.808 2.913 0.858 ;
      RECT 2.863 0.858 2.913 1.166 ;
      RECT 2.823 0.354 2.873 0.808 ;
      RECT 1.747 0.88 1.949 0.93 ;
      RECT 1.747 0.673 2.093 0.723 ;
      RECT 1.607 1.317 1.949 1.367 ;
      RECT 1.607 1.367 1.657 1.528 ;
      RECT 1.403 1.528 1.657 1.578 ;
      RECT 1.747 0.723 1.797 0.88 ;
      RECT 1.899 0.93 1.949 1.317 ;
      RECT 0.947 0.626 1.333 0.676 ;
      RECT 1.039 0.676 1.089 1.152 ;
      RECT 1.039 0.401 1.089 0.626 ;
      RECT 0.548 0.573 0.725 0.623 ;
      RECT 0.279 0.844 0.598 0.894 ;
      RECT 0.548 0.623 0.598 0.844 ;
      RECT 0.279 0.601 0.369 0.651 ;
      RECT 0.279 0.455 0.329 0.601 ;
      RECT 0.319 0.651 0.369 0.844 ;
      RECT 0.279 0.894 0.329 1.246 ;
      RECT 2.771 1.528 3.461 1.578 ;
      RECT 3.227 0.577 3.578 0.627 ;
      RECT 3.528 0.704 4.034 0.754 ;
      RECT 3.984 0.654 4.034 0.704 ;
      RECT 3.984 0.604 4.221 0.654 ;
      RECT 3.528 0.754 3.578 0.758 ;
      RECT 3.528 0.627 3.578 0.704 ;
      RECT 0.567 0.301 0.953 0.351 ;
      RECT 0.583 1.316 0.954 1.366 ;
      RECT 0.583 0.98 0.633 1.316 ;
      RECT 0.947 0.104 1.789 0.154 ;
      RECT 1.571 0.154 1.621 0.217 ;
      RECT 1.707 1.417 2.093 1.467 ;
    LAYER PO ;
      RECT 2.037 0.966 2.067 1.606 ;
      RECT 1.125 0.076 1.155 1.606 ;
      RECT 2.189 0.076 2.219 1.606 ;
      RECT 0.669 0.87 0.699 1.606 ;
      RECT 1.581 0.076 1.611 0.597 ;
      RECT 2.645 1.032 2.675 1.606 ;
      RECT 0.365 0.076 0.395 1.606 ;
      RECT 3.405 0.076 3.435 0.755 ;
      RECT 3.557 0.076 3.587 1.606 ;
      RECT 0.669 0.076 0.699 0.651 ;
      RECT 4.469 0.076 4.499 1.606 ;
      RECT 1.581 0.92 1.611 1.606 ;
      RECT 3.709 0.076 3.739 1.606 ;
      RECT 1.429 0.076 1.459 1.606 ;
      RECT 4.165 0.076 4.195 1.606 ;
      RECT 4.013 0.076 4.043 1.606 ;
      RECT 4.317 0.076 4.347 1.606 ;
      RECT 3.861 0.076 3.891 1.606 ;
      RECT 1.885 0.076 1.915 1.606 ;
      RECT 1.277 0.076 1.307 1.606 ;
      RECT 2.341 0.076 2.371 1.606 ;
      RECT 3.405 1.132 3.435 1.606 ;
      RECT 2.037 0.076 2.067 0.751 ;
      RECT 2.949 0.076 2.979 1.606 ;
      RECT 3.253 0.076 3.283 1.606 ;
      RECT 1.733 0.076 1.763 1.606 ;
      RECT 3.101 0.076 3.131 1.606 ;
      RECT 0.973 0.076 1.003 1.606 ;
      RECT 2.645 0.076 2.675 0.597 ;
      RECT 2.493 0.076 2.523 1.606 ;
      RECT 0.517 0.076 0.547 0.597 ;
      RECT 0.517 0.816 0.547 1.606 ;
      RECT 2.797 0.076 2.827 1.606 ;
      RECT 0.821 0.076 0.851 1.606 ;
      RECT 0.061 0.076 0.091 1.606 ;
      RECT 0.213 0.076 0.243 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 4.675 1.773 ;
  END
END DFFSSRX2_RVT

MACRO NAND3X0_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.064 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.739 0.705 0.781 ;
      LAYER M1 ;
        RECT 0.705 0.785 0.815 0.815 ;
        RECT 0.643 0.735 0.815 0.785 ;
        RECT 0.705 0.705 0.815 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.891 0.553 0.933 ;
      LAYER M1 ;
        RECT 0.553 0.937 0.663 0.967 ;
        RECT 0.491 0.887 0.663 0.937 ;
        RECT 0.553 0.857 0.663 0.887 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.891 0.401 0.933 ;
      LAYER M1 ;
        RECT 0.249 0.937 0.359 0.967 ;
        RECT 0.249 0.887 0.421 0.937 ;
        RECT 0.249 0.857 0.359 0.887 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END A3
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.739 0.141 0.781 0.183 ;
        RECT 0.739 0.233 0.781 0.275 ;
        RECT 0.739 0.325 0.781 0.367 ;
        RECT 0.739 0.417 0.781 0.459 ;
        RECT 0.435 1.213 0.477 1.255 ;
        RECT 0.739 1.213 0.781 1.255 ;
        RECT 0.435 1.305 0.477 1.347 ;
        RECT 0.739 1.305 0.781 1.347 ;
        RECT 0.435 1.397 0.477 1.439 ;
        RECT 0.739 1.397 0.781 1.439 ;
        RECT 0.435 1.489 0.477 1.531 ;
        RECT 0.739 1.489 0.781 1.531 ;
      LAYER M1 ;
        RECT 0.431 1.14 0.481 1.551 ;
        RECT 0.735 1.14 0.785 1.551 ;
        RECT 0.431 1.091 0.915 1.14 ;
        RECT 0.456 1.09 0.915 1.091 ;
        RECT 0.865 0.967 0.915 1.09 ;
        RECT 0.855 0.857 0.967 0.967 ;
        RECT 0.865 0.655 0.915 0.857 ;
        RECT 0.735 0.605 0.915 0.655 ;
        RECT 0.735 0.106 0.785 0.605 ;
    END
    ANTENNADIFFAREA 0.1348 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.213 0.325 1.255 ;
        RECT 0.587 1.213 0.629 1.255 ;
        RECT 0.283 1.305 0.325 1.347 ;
        RECT 0.587 1.305 0.629 1.347 ;
        RECT 0.283 1.397 0.325 1.439 ;
        RECT 0.587 1.397 0.629 1.439 ;
        RECT 0.283 1.489 0.325 1.531 ;
        RECT 0.587 1.489 0.629 1.531 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.064 1.702 ;
        RECT 0.279 1.193 0.329 1.642 ;
        RECT 0.583 1.193 0.633 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 0.283 0.141 0.325 0.183 ;
        RECT 0.283 0.233 0.325 0.275 ;
        RECT 0.283 0.325 0.325 0.367 ;
        RECT 0.283 0.417 0.325 0.459 ;
      LAYER M1 ;
        RECT 0.279 0.03 0.329 0.479 ;
        RECT 0 -0.03 1.064 0.03 ;
    END
  END VSS
  OBS
    LAYER PO ;
      RECT 0.061 0.071 0.091 1.61 ;
      RECT 0.821 0.071 0.851 1.61 ;
      RECT 0.213 0.071 0.243 1.61 ;
      RECT 0.517 0.071 0.547 1.61 ;
      RECT 0.365 0.071 0.395 1.61 ;
      RECT 0.669 0.071 0.699 1.61 ;
      RECT 0.973 0.071 1.003 1.61 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.178 1.773 ;
  END
END NAND3X0_RVT

MACRO AND2X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.368 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.887 0.553 0.929 ;
      LAYER M1 ;
        RECT 0.401 0.933 0.511 0.967 ;
        RECT 0.401 0.883 0.573 0.933 ;
        RECT 0.401 0.857 0.511 0.883 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.249 0.785 0.359 0.815 ;
        RECT 0.249 0.735 0.421 0.785 ;
        RECT 0.249 0.705 0.359 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.739 0.15 0.781 0.192 ;
        RECT 1.043 0.15 1.085 0.192 ;
        RECT 0.739 0.242 0.781 0.284 ;
        RECT 1.043 0.242 1.085 0.284 ;
        RECT 0.739 0.334 0.781 0.376 ;
        RECT 1.043 0.334 1.085 0.376 ;
        RECT 0.739 0.426 0.781 0.468 ;
        RECT 1.043 0.426 1.085 0.468 ;
        RECT 0.739 0.838 0.781 0.88 ;
        RECT 1.043 0.838 1.085 0.88 ;
        RECT 0.739 0.93 0.781 0.972 ;
        RECT 1.043 0.93 1.085 0.972 ;
        RECT 0.739 1.022 0.781 1.064 ;
        RECT 1.043 1.022 1.085 1.064 ;
        RECT 0.739 1.114 0.781 1.156 ;
        RECT 1.043 1.114 1.085 1.156 ;
        RECT 0.739 1.206 0.781 1.248 ;
        RECT 1.043 1.206 1.085 1.248 ;
        RECT 0.739 1.298 0.781 1.34 ;
        RECT 1.043 1.298 1.085 1.34 ;
        RECT 0.739 1.39 0.781 1.432 ;
        RECT 1.043 1.39 1.085 1.432 ;
        RECT 0.739 1.482 0.781 1.524 ;
        RECT 1.043 1.482 1.085 1.524 ;
      LAYER M1 ;
        RECT 0.735 0.753 0.785 1.544 ;
        RECT 1.039 0.753 1.089 1.544 ;
        RECT 0.735 0.703 1.181 0.753 ;
        RECT 1.131 0.663 1.181 0.703 ;
        RECT 1.131 0.553 1.271 0.663 ;
        RECT 0.735 0.503 1.181 0.553 ;
        RECT 0.735 0.13 0.785 0.503 ;
        RECT 1.039 0.13 1.089 0.503 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.891 0.838 0.933 0.88 ;
        RECT 0.891 0.93 0.933 0.972 ;
        RECT 0.891 1.022 0.933 1.064 ;
        RECT 0.891 1.114 0.933 1.156 ;
        RECT 0.891 1.206 0.933 1.248 ;
        RECT 0.435 1.215 0.477 1.257 ;
        RECT 0.891 1.298 0.933 1.34 ;
        RECT 0.435 1.307 0.477 1.349 ;
        RECT 0.891 1.39 0.933 1.432 ;
        RECT 0.435 1.399 0.477 1.441 ;
        RECT 0.891 1.482 0.933 1.524 ;
        RECT 0.435 1.491 0.477 1.533 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.368 1.702 ;
        RECT 0.431 1.195 0.481 1.642 ;
        RECT 0.887 0.818 0.937 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 0.283 0.141 0.325 0.183 ;
        RECT 0.891 0.152 0.933 0.194 ;
        RECT 0.283 0.233 0.325 0.275 ;
        RECT 0.891 0.244 0.933 0.286 ;
        RECT 0.283 0.325 0.325 0.367 ;
        RECT 0.891 0.336 0.933 0.378 ;
        RECT 0.283 0.417 0.325 0.459 ;
      LAYER M1 ;
        RECT 0.279 0.03 0.329 0.479 ;
        RECT 0.887 0.03 0.937 0.398 ;
        RECT 0 -0.03 1.368 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.149 0.603 1.029 0.653 ;
      RECT 0.149 0.608 0.199 1.079 ;
      RECT 0.279 1.029 0.329 1.553 ;
      RECT 0.15 1.029 0.633 1.079 ;
      RECT 0.583 1.053 0.633 1.553 ;
      RECT 0.583 0.121 0.633 0.647 ;
    LAYER PO ;
      RECT 0.973 0.072 1.003 1.604 ;
      RECT 1.125 0.072 1.155 1.603 ;
      RECT 0.821 0.072 0.851 1.604 ;
      RECT 0.669 0.071 0.699 1.603 ;
      RECT 0.365 0.071 0.395 1.603 ;
      RECT 0.517 0.071 0.547 1.603 ;
      RECT 0.213 0.071 0.243 1.603 ;
      RECT 0.061 0.071 0.091 1.603 ;
      RECT 1.277 0.072 1.307 1.61 ;
    LAYER CO ;
      RECT 0.587 0.417 0.629 0.459 ;
      RECT 0.587 1.491 0.629 1.533 ;
      RECT 0.587 1.399 0.629 1.441 ;
      RECT 0.815 0.607 0.857 0.649 ;
      RECT 0.587 0.233 0.629 0.275 ;
      RECT 0.587 0.141 0.629 0.183 ;
      RECT 0.967 0.607 1.009 0.649 ;
      RECT 0.587 1.215 0.629 1.257 ;
      RECT 0.587 1.307 0.629 1.349 ;
      RECT 0.283 1.215 0.325 1.257 ;
      RECT 0.283 1.307 0.325 1.349 ;
      RECT 0.283 1.491 0.325 1.533 ;
      RECT 0.283 1.399 0.325 1.441 ;
      RECT 0.587 0.325 0.629 0.367 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.483 1.773 ;
  END
END AND2X2_RVT

MACRO INVX0_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.684 0.401 0.726 ;
      LAYER M1 ;
        RECT 0.249 0.73 0.362 0.815 ;
        RECT 0.249 0.68 0.421 0.73 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.435 0.325 0.477 0.367 ;
        RECT 0.435 0.417 0.477 0.459 ;
        RECT 0.435 0.509 0.477 0.551 ;
        RECT 0.435 0.843 0.477 0.885 ;
        RECT 0.435 0.935 0.477 0.977 ;
        RECT 0.435 1.027 0.477 1.069 ;
        RECT 0.435 1.119 0.477 1.161 ;
        RECT 0.435 1.211 0.477 1.253 ;
      LAYER M1 ;
        RECT 0.431 0.873 0.481 1.288 ;
        RECT 0.431 0.823 0.521 0.873 ;
        RECT 0.471 0.663 0.521 0.823 ;
        RECT 0.471 0.587 0.663 0.663 ;
        RECT 0.431 0.537 0.663 0.587 ;
        RECT 0.431 0.305 0.481 0.537 ;
    END
    ANTENNADIFFAREA 0.0805 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 0.948 0.325 0.99 ;
        RECT 0.283 1.04 0.325 1.082 ;
        RECT 0.283 1.132 0.325 1.174 ;
        RECT 0.283 1.224 0.325 1.266 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 0.76 1.702 ;
        RECT 0.279 0.928 0.329 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.283 0.318 0.325 0.36 ;
        RECT 0.283 0.41 0.325 0.452 ;
        RECT 0.283 0.502 0.325 0.544 ;
      LAYER M1 ;
        RECT 0.279 0.03 0.329 0.564 ;
        RECT 0 -0.03 0.76 0.03 ;
    END
  END VSS
  OBS
    LAYER PO ;
      RECT 0.213 0.071 0.243 1.606 ;
      RECT 0.365 0.069 0.395 1.606 ;
      RECT 0.669 0.071 0.699 1.606 ;
      RECT 0.517 0.071 0.547 1.606 ;
      RECT 0.061 0.071 0.091 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 0.875 1.773 ;
  END
END INVX0_RVT

MACRO AND3X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.739 0.705 0.781 ;
      LAYER M1 ;
        RECT 0.553 0.785 0.663 0.815 ;
        RECT 0.553 0.735 0.725 0.785 ;
        RECT 0.553 0.705 0.663 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.043 0.553 1.085 ;
      LAYER M1 ;
        RECT 0.401 1.089 0.511 1.119 ;
        RECT 0.401 1.039 0.573 1.089 ;
        RECT 0.401 1.009 0.511 1.039 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.249 0.785 0.359 0.815 ;
        RECT 0.249 0.735 0.421 0.785 ;
        RECT 0.249 0.705 0.359 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END A3
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.891 0.149 0.933 0.191 ;
        RECT 1.195 0.149 1.237 0.191 ;
        RECT 0.891 0.241 0.933 0.283 ;
        RECT 1.195 0.241 1.237 0.283 ;
        RECT 0.891 0.333 0.933 0.375 ;
        RECT 1.195 0.333 1.237 0.375 ;
        RECT 0.891 0.425 0.933 0.467 ;
        RECT 1.195 0.425 1.237 0.467 ;
        RECT 0.891 0.838 0.933 0.88 ;
        RECT 1.195 0.838 1.237 0.88 ;
        RECT 0.891 0.93 0.933 0.972 ;
        RECT 1.195 0.93 1.237 0.972 ;
        RECT 0.891 1.022 0.933 1.064 ;
        RECT 1.195 1.022 1.237 1.064 ;
        RECT 0.891 1.114 0.933 1.156 ;
        RECT 1.195 1.114 1.237 1.156 ;
        RECT 0.891 1.206 0.933 1.248 ;
        RECT 1.195 1.206 1.237 1.248 ;
        RECT 0.891 1.298 0.933 1.34 ;
        RECT 1.195 1.298 1.237 1.34 ;
        RECT 0.891 1.39 0.933 1.432 ;
        RECT 1.195 1.39 1.237 1.432 ;
        RECT 0.891 1.482 0.933 1.524 ;
        RECT 1.195 1.482 1.237 1.524 ;
      LAYER M1 ;
        RECT 0.887 0.764 0.937 1.544 ;
        RECT 1.191 0.764 1.241 1.544 ;
        RECT 0.887 0.714 1.328 0.764 ;
        RECT 1.278 0.663 1.328 0.714 ;
        RECT 1.278 0.553 1.423 0.663 ;
        RECT 1.278 0.529 1.328 0.553 ;
        RECT 0.887 0.479 1.328 0.529 ;
        RECT 0.887 0.129 0.937 0.479 ;
        RECT 1.191 0.129 1.241 0.479 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.043 0.838 1.085 0.88 ;
        RECT 1.043 0.93 1.085 0.972 ;
        RECT 1.043 1.022 1.085 1.064 ;
        RECT 1.043 1.114 1.085 1.156 ;
        RECT 1.043 1.206 1.085 1.248 ;
        RECT 1.043 1.298 1.085 1.34 ;
        RECT 1.043 1.39 1.085 1.432 ;
        RECT 0.283 1.399 0.325 1.441 ;
        RECT 0.587 1.399 0.629 1.441 ;
        RECT 1.043 1.482 1.085 1.524 ;
        RECT 0.283 1.491 0.325 1.533 ;
        RECT 0.587 1.491 0.629 1.533 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.52 1.702 ;
        RECT 0.279 1.379 0.329 1.642 ;
        RECT 0.583 1.379 0.633 1.642 ;
        RECT 1.039 0.814 1.089 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 0.283 0.141 0.325 0.183 ;
        RECT 1.043 0.151 1.085 0.193 ;
        RECT 0.283 0.233 0.325 0.275 ;
        RECT 1.043 0.243 1.085 0.285 ;
        RECT 0.283 0.325 0.325 0.367 ;
        RECT 1.043 0.335 1.085 0.377 ;
        RECT 0.283 0.417 0.325 0.459 ;
      LAYER M1 ;
        RECT 0.279 0.03 0.329 0.479 ;
        RECT 1.041 0.03 1.091 0.398 ;
        RECT 0 -0.03 1.52 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.735 0.614 1.181 0.664 ;
      RECT 0.431 1.187 0.481 1.553 ;
      RECT 0.735 1.187 0.785 1.553 ;
      RECT 0.456 1.187 0.825 1.237 ;
      RECT 0.775 0.614 0.825 1.211 ;
      RECT 0.735 0.121 0.785 0.642 ;
    LAYER PO ;
      RECT 1.125 0.071 1.155 1.604 ;
      RECT 1.277 0.072 1.307 1.603 ;
      RECT 0.973 0.071 1.003 1.604 ;
      RECT 1.429 0.072 1.459 1.603 ;
      RECT 0.669 0.071 0.699 1.603 ;
      RECT 0.365 0.071 0.395 1.603 ;
      RECT 0.517 0.071 0.547 1.603 ;
      RECT 0.213 0.071 0.243 1.603 ;
      RECT 0.821 0.071 0.851 1.603 ;
      RECT 0.061 0.071 0.091 1.603 ;
    LAYER CO ;
      RECT 1.119 0.618 1.161 0.66 ;
      RECT 0.967 0.618 1.009 0.66 ;
      RECT 0.435 1.491 0.477 1.533 ;
      RECT 0.435 1.399 0.477 1.441 ;
      RECT 0.739 1.399 0.781 1.441 ;
      RECT 0.739 0.141 0.781 0.183 ;
      RECT 0.739 0.233 0.781 0.275 ;
      RECT 0.739 0.325 0.781 0.367 ;
      RECT 0.739 0.417 0.781 0.459 ;
      RECT 0.739 1.491 0.781 1.533 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.635 1.773 ;
  END
END AND3X2_RVT

MACRO AND4X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 1.043 0.857 1.085 ;
      LAYER M1 ;
        RECT 0.705 1.089 0.815 1.119 ;
        RECT 0.705 1.039 0.877 1.089 ;
        RECT 0.705 1.009 0.815 1.039 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0183 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.739 0.705 0.781 ;
      LAYER M1 ;
        RECT 0.553 0.785 0.663 0.815 ;
        RECT 0.553 0.735 0.725 0.785 ;
        RECT 0.553 0.705 0.663 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0183 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.043 0.553 1.085 ;
      LAYER M1 ;
        RECT 0.401 1.089 0.511 1.119 ;
        RECT 0.401 1.039 0.573 1.089 ;
        RECT 0.401 1.009 0.511 1.039 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0183 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.249 0.785 0.359 0.815 ;
        RECT 0.249 0.735 0.421 0.785 ;
        RECT 0.249 0.705 0.359 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0183 ;
  END A4
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.195 0.15 1.237 0.192 ;
        RECT 1.195 0.242 1.237 0.284 ;
        RECT 1.195 0.334 1.237 0.376 ;
        RECT 1.195 0.426 1.237 0.468 ;
        RECT 1.195 0.851 1.237 0.893 ;
        RECT 1.195 0.943 1.237 0.985 ;
        RECT 1.195 1.035 1.237 1.077 ;
        RECT 1.195 1.127 1.237 1.169 ;
        RECT 1.195 1.219 1.237 1.261 ;
        RECT 1.195 1.311 1.237 1.353 ;
        RECT 1.195 1.403 1.237 1.445 ;
        RECT 1.195 1.495 1.237 1.537 ;
      LAYER M1 ;
        RECT 1.191 0.805 1.241 1.557 ;
        RECT 1.191 0.755 1.34 0.805 ;
        RECT 1.29 0.663 1.34 0.755 ;
        RECT 1.29 0.601 1.423 0.663 ;
        RECT 1.191 0.553 1.423 0.601 ;
        RECT 1.191 0.551 1.315 0.553 ;
        RECT 1.191 0.117 1.241 0.551 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.043 0.851 1.085 0.893 ;
        RECT 1.043 0.943 1.085 0.985 ;
        RECT 1.043 1.035 1.085 1.077 ;
        RECT 1.043 1.127 1.085 1.169 ;
        RECT 1.043 1.219 1.085 1.261 ;
        RECT 1.043 1.311 1.085 1.353 ;
        RECT 1.043 1.403 1.085 1.445 ;
        RECT 0.435 1.405 0.477 1.447 ;
        RECT 0.739 1.405 0.781 1.447 ;
        RECT 1.043 1.495 1.085 1.537 ;
        RECT 0.435 1.497 0.477 1.539 ;
        RECT 0.739 1.497 0.781 1.539 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.52 1.702 ;
        RECT 0.431 1.385 0.481 1.642 ;
        RECT 0.735 1.385 0.785 1.642 ;
        RECT 1.039 0.831 1.089 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 0.283 0.141 0.325 0.183 ;
        RECT 1.043 0.15 1.085 0.192 ;
        RECT 0.283 0.233 0.325 0.275 ;
        RECT 1.043 0.242 1.085 0.284 ;
        RECT 0.283 0.325 0.325 0.367 ;
        RECT 1.043 0.334 1.085 0.376 ;
        RECT 0.283 0.417 0.325 0.459 ;
        RECT 1.043 0.426 1.085 0.468 ;
      LAYER M1 ;
        RECT 1.039 0.03 1.089 0.488 ;
        RECT 0.279 0.03 0.329 0.479 ;
        RECT 0 -0.03 1.52 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.97 0.656 1.181 0.706 ;
      RECT 0.279 1.263 0.329 1.559 ;
      RECT 0.583 1.289 0.633 1.559 ;
      RECT 0.927 0.622 0.977 1.288 ;
      RECT 0.887 0.622 0.97 0.672 ;
      RECT 0.887 0.121 0.937 0.647 ;
      RECT 0.279 1.263 0.977 1.313 ;
      RECT 0.887 1.279 0.937 1.559 ;
    LAYER PO ;
      RECT 1.277 0.072 1.307 1.609 ;
      RECT 1.429 0.072 1.459 1.609 ;
      RECT 1.125 0.072 1.155 1.609 ;
      RECT 0.973 0.071 1.003 1.609 ;
      RECT 0.669 0.071 0.699 1.609 ;
      RECT 0.365 0.071 0.395 1.609 ;
      RECT 0.517 0.071 0.547 1.609 ;
      RECT 0.213 0.071 0.243 1.609 ;
      RECT 0.821 0.071 0.851 1.609 ;
      RECT 0.061 0.071 0.091 1.609 ;
    LAYER CO ;
      RECT 0.891 0.417 0.933 0.459 ;
      RECT 0.891 0.325 0.933 0.367 ;
      RECT 0.891 0.233 0.933 0.275 ;
      RECT 0.891 0.141 0.933 0.183 ;
      RECT 1.119 0.66 1.161 0.702 ;
      RECT 0.891 1.405 0.933 1.447 ;
      RECT 0.891 1.497 0.933 1.539 ;
      RECT 0.283 1.405 0.325 1.447 ;
      RECT 0.283 1.497 0.325 1.539 ;
      RECT 0.587 1.405 0.629 1.447 ;
      RECT 0.587 1.497 0.629 1.539 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.635 1.773 ;
  END
END AND4X1_RVT

MACRO OA22X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.271 0.81 0.421 0.817 ;
        RECT 0.249 0.71 0.421 0.81 ;
        RECT 0.249 0.701 0.359 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0216 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.482 0.553 1.524 ;
      LAYER M1 ;
        RECT 0.401 1.571 0.511 1.575 ;
        RECT 0.401 1.464 0.573 1.571 ;
        RECT 0.426 1.46 0.573 1.464 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0216 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.744 0.857 0.786 ;
      LAYER M1 ;
        RECT 0.811 1.002 0.968 1.139 ;
        RECT 0.811 0.715 0.861 1.002 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0216 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.747 0.705 0.789 ;
      LAYER M1 ;
        RECT 0.56 0.963 0.709 0.986 ;
        RECT 0.553 0.854 0.709 0.963 ;
        RECT 0.659 0.723 0.709 0.854 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0216 ;
  END A4
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.195 0.239 1.237 0.281 ;
        RECT 1.195 0.331 1.237 0.373 ;
        RECT 1.195 0.423 1.237 0.465 ;
        RECT 1.195 0.987 1.237 1.029 ;
        RECT 1.195 1.079 1.237 1.121 ;
        RECT 1.195 1.171 1.237 1.213 ;
        RECT 1.195 1.263 1.237 1.305 ;
        RECT 1.195 1.355 1.237 1.397 ;
      LAYER M1 ;
        RECT 1.191 1.006 1.241 1.426 ;
        RECT 1.191 0.956 1.38 1.006 ;
        RECT 1.33 0.542 1.38 0.956 ;
        RECT 1.191 0.53 1.38 0.542 ;
        RECT 1.191 0.492 1.455 0.53 ;
        RECT 1.191 0.188 1.241 0.492 ;
        RECT 1.295 0.392 1.455 0.492 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.079 0.325 1.121 ;
        RECT 0.283 1.171 0.325 1.213 ;
        RECT 0.283 1.263 0.325 1.305 ;
        RECT 0.283 1.355 0.325 1.397 ;
        RECT 0.891 1.355 0.933 1.397 ;
        RECT 1.043 1.355 1.085 1.397 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.52 1.702 ;
        RECT 0.279 0.958 0.329 1.642 ;
        RECT 0.887 1.335 0.937 1.642 ;
        RECT 1.039 1.333 1.089 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.043 0.203 1.085 0.245 ;
        RECT 0.435 0.239 0.477 0.281 ;
        RECT 1.043 0.295 1.085 0.337 ;
        RECT 0.435 0.331 0.477 0.373 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.512 ;
        RECT 1.039 0.03 1.089 0.399 ;
        RECT 0 -0.03 1.52 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.079 0.699 1.129 1.226 ;
      RECT 0.735 0.613 1.165 0.663 ;
      RECT 1.079 0.663 1.165 0.699 ;
      RECT 0.583 1.226 1.129 1.276 ;
      RECT 0.735 0.212 0.785 0.613 ;
      RECT 0.583 1.276 0.633 1.393 ;
      RECT 0.583 1.106 0.633 1.226 ;
      RECT 0.583 0.095 0.937 0.145 ;
      RECT 0.279 0.598 0.633 0.648 ;
      RECT 0.583 0.145 0.633 0.598 ;
      RECT 0.887 0.145 0.937 0.504 ;
      RECT 0.279 0.178 0.329 0.598 ;
    LAYER PO ;
      RECT 0.061 0.101 0.091 1.469 ;
      RECT 0.517 0.101 0.547 1.567 ;
      RECT 0.213 0.101 0.243 1.469 ;
      RECT 0.973 0.101 1.003 1.469 ;
      RECT 0.821 0.101 0.851 1.469 ;
      RECT 0.669 0.101 0.699 1.469 ;
      RECT 1.125 0.069 1.155 1.608 ;
      RECT 0.365 0.101 0.395 1.469 ;
      RECT 1.277 0.101 1.307 1.469 ;
      RECT 1.429 0.101 1.459 1.469 ;
    LAYER CO ;
      RECT 0.891 0.331 0.933 0.373 ;
      RECT 0.891 0.239 0.933 0.281 ;
      RECT 0.739 0.331 0.781 0.373 ;
      RECT 0.283 0.331 0.325 0.373 ;
      RECT 0.739 0.239 0.781 0.281 ;
      RECT 0.283 0.239 0.325 0.281 ;
      RECT 0.587 0.331 0.629 0.373 ;
      RECT 0.587 0.239 0.629 0.281 ;
      RECT 1.119 0.635 1.161 0.677 ;
      RECT 0.587 1.23 0.629 1.272 ;
      RECT 0.587 1.138 0.629 1.18 ;
      RECT 0.587 1.322 0.629 1.364 ;
    LAYER NWELL ;
      RECT -0.135 0.679 1.636 1.787 ;
  END
END OA22X1_RVT

MACRO INVX2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.912 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.664 0.401 0.706 ;
        RECT 0.511 0.664 0.553 0.706 ;
      LAYER M1 ;
        RECT 0.249 0.71 0.362 0.815 ;
        RECT 0.249 0.66 0.588 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0732 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.283 0.151 0.325 0.193 ;
        RECT 0.587 0.151 0.629 0.193 ;
        RECT 0.283 0.243 0.325 0.285 ;
        RECT 0.587 0.243 0.629 0.285 ;
        RECT 0.283 0.335 0.325 0.377 ;
        RECT 0.587 0.335 0.629 0.377 ;
        RECT 0.283 0.427 0.325 0.469 ;
        RECT 0.587 0.427 0.629 0.469 ;
        RECT 0.283 1.027 0.325 1.069 ;
        RECT 0.587 1.027 0.629 1.069 ;
        RECT 0.283 1.119 0.325 1.161 ;
        RECT 0.587 1.119 0.629 1.161 ;
        RECT 0.283 1.211 0.325 1.253 ;
        RECT 0.587 1.211 0.629 1.253 ;
        RECT 0.283 1.303 0.325 1.345 ;
        RECT 0.587 1.303 0.629 1.345 ;
        RECT 0.283 1.395 0.325 1.437 ;
        RECT 0.587 1.395 0.629 1.437 ;
        RECT 0.283 1.487 0.325 1.529 ;
        RECT 0.587 1.487 0.629 1.529 ;
      LAYER M1 ;
        RECT 0.279 0.942 0.329 1.564 ;
        RECT 0.583 0.942 0.633 1.564 ;
        RECT 0.279 0.892 0.689 0.942 ;
        RECT 0.639 0.663 0.689 0.892 ;
        RECT 0.639 0.587 0.815 0.663 ;
        RECT 0.279 0.537 0.815 0.587 ;
        RECT 0.279 0.116 0.329 0.537 ;
        RECT 0.583 0.116 0.633 0.537 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.435 1.027 0.477 1.069 ;
        RECT 0.435 1.119 0.477 1.161 ;
        RECT 0.435 1.211 0.477 1.253 ;
        RECT 0.435 1.303 0.477 1.345 ;
        RECT 0.435 1.395 0.477 1.437 ;
        RECT 0.435 1.487 0.477 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 0.912 1.702 ;
        RECT 0.431 0.992 0.481 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.435 0.149 0.477 0.191 ;
        RECT 0.435 0.241 0.477 0.283 ;
        RECT 0.435 0.333 0.477 0.375 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.41 ;
        RECT 0 -0.03 0.912 0.03 ;
    END
  END VSS
  OBS
    LAYER PO ;
      RECT 0.213 0.071 0.243 1.606 ;
      RECT 0.365 0.069 0.395 1.606 ;
      RECT 0.821 0.071 0.851 1.606 ;
      RECT 0.669 0.071 0.699 1.606 ;
      RECT 0.517 0.069 0.547 1.606 ;
      RECT 0.061 0.071 0.091 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.027 1.773 ;
  END
END INVX2_RVT

MACRO NBUFFX4_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.659 0.401 0.701 ;
      LAYER M1 ;
        RECT 0.249 0.705 0.362 0.815 ;
        RECT 0.249 0.655 0.436 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.587 0.151 0.629 0.193 ;
        RECT 0.891 0.151 0.933 0.193 ;
        RECT 1.195 0.151 1.237 0.193 ;
        RECT 0.587 0.243 0.629 0.285 ;
        RECT 0.891 0.243 0.933 0.285 ;
        RECT 1.195 0.243 1.237 0.285 ;
        RECT 0.587 0.335 0.629 0.377 ;
        RECT 0.891 0.335 0.933 0.377 ;
        RECT 1.195 0.335 1.237 0.377 ;
        RECT 0.587 0.427 0.629 0.469 ;
        RECT 0.891 0.427 0.933 0.469 ;
        RECT 1.195 0.427 1.237 0.469 ;
        RECT 0.587 1.027 0.629 1.069 ;
        RECT 0.891 1.027 0.933 1.069 ;
        RECT 1.195 1.027 1.237 1.069 ;
        RECT 0.587 1.119 0.629 1.161 ;
        RECT 0.891 1.119 0.933 1.161 ;
        RECT 1.195 1.119 1.237 1.161 ;
        RECT 0.587 1.211 0.629 1.253 ;
        RECT 0.891 1.211 0.933 1.253 ;
        RECT 1.195 1.211 1.237 1.253 ;
        RECT 0.587 1.303 0.629 1.345 ;
        RECT 0.891 1.303 0.933 1.345 ;
        RECT 1.195 1.303 1.237 1.345 ;
        RECT 0.587 1.395 0.629 1.437 ;
        RECT 0.891 1.395 0.933 1.437 ;
        RECT 1.195 1.395 1.237 1.437 ;
        RECT 0.587 1.487 0.629 1.529 ;
        RECT 0.891 1.487 0.933 1.529 ;
        RECT 1.195 1.487 1.237 1.529 ;
      LAYER M1 ;
        RECT 0.583 0.942 0.633 1.564 ;
        RECT 0.887 0.942 0.937 1.564 ;
        RECT 1.191 0.942 1.241 1.564 ;
        RECT 0.583 0.892 1.296 0.942 ;
        RECT 1.246 0.663 1.296 0.892 ;
        RECT 1.246 0.587 1.423 0.663 ;
        RECT 0.583 0.537 1.423 0.587 ;
        RECT 0.583 0.116 0.633 0.537 ;
        RECT 0.887 0.116 0.937 0.537 ;
        RECT 1.191 0.116 1.241 0.537 ;
    END
    ANTENNADIFFAREA 0.3976 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.022 0.325 1.064 ;
        RECT 0.739 1.027 0.781 1.069 ;
        RECT 1.043 1.027 1.085 1.069 ;
        RECT 0.283 1.114 0.325 1.156 ;
        RECT 0.739 1.119 0.781 1.161 ;
        RECT 1.043 1.119 1.085 1.161 ;
        RECT 0.283 1.206 0.325 1.248 ;
        RECT 0.739 1.211 0.781 1.253 ;
        RECT 1.043 1.211 1.085 1.253 ;
        RECT 0.283 1.298 0.325 1.34 ;
        RECT 0.739 1.303 0.781 1.345 ;
        RECT 1.043 1.303 1.085 1.345 ;
        RECT 0.283 1.39 0.325 1.432 ;
        RECT 0.739 1.395 0.781 1.437 ;
        RECT 1.043 1.395 1.085 1.437 ;
        RECT 0.283 1.482 0.325 1.524 ;
        RECT 0.739 1.487 0.781 1.529 ;
        RECT 1.043 1.487 1.085 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.52 1.702 ;
        RECT 0.279 0.987 0.329 1.642 ;
        RECT 0.735 0.992 0.785 1.642 ;
        RECT 1.039 0.992 1.089 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 0.283 0.144 0.325 0.186 ;
        RECT 0.739 0.149 0.781 0.191 ;
        RECT 1.043 0.149 1.085 0.191 ;
        RECT 0.283 0.236 0.325 0.278 ;
        RECT 0.739 0.241 0.781 0.283 ;
        RECT 1.043 0.241 1.085 0.283 ;
        RECT 0.283 0.328 0.325 0.37 ;
        RECT 0.739 0.333 0.781 0.375 ;
        RECT 1.043 0.333 1.085 0.375 ;
      LAYER M1 ;
        RECT 0.735 0.03 0.785 0.41 ;
        RECT 1.039 0.03 1.089 0.41 ;
        RECT 0.279 0.03 0.329 0.405 ;
        RECT 0 -0.03 1.52 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.435 1.022 0.477 1.064 ;
      RECT 0.435 1.114 0.477 1.156 ;
      RECT 0.435 1.022 0.477 1.064 ;
      RECT 0.435 1.482 0.477 1.524 ;
      RECT 0.435 1.482 0.477 1.524 ;
      RECT 0.435 1.39 0.477 1.432 ;
      RECT 0.435 0.146 0.477 0.188 ;
      RECT 0.435 0.238 0.477 0.28 ;
      RECT 0.435 0.33 0.477 0.372 ;
      RECT 0.435 0.33 0.477 0.372 ;
      RECT 0.435 0.422 0.477 0.464 ;
      RECT 1.119 0.664 1.161 0.706 ;
      RECT 0.967 0.664 1.009 0.706 ;
      RECT 0.435 0.146 0.477 0.188 ;
      RECT 0.435 1.298 0.477 1.34 ;
      RECT 0.435 1.298 0.477 1.34 ;
      RECT 0.435 1.206 0.477 1.248 ;
      RECT 0.663 0.664 0.705 0.706 ;
      RECT 0.815 0.664 0.857 0.706 ;
      RECT 0.435 1.206 0.477 1.248 ;
      RECT 0.435 1.39 0.477 1.432 ;
      RECT 0.435 1.114 0.477 1.156 ;
    LAYER M1 ;
      RECT 0.487 0.66 1.196 0.71 ;
      RECT 0.456 0.822 0.537 0.872 ;
      RECT 0.487 0.609 0.537 0.872 ;
      RECT 0.431 0.822 0.481 1.559 ;
      RECT 0.483 0.532 0.533 0.637 ;
      RECT 0.431 0.887 0.474 0.937 ;
      RECT 0.431 0.532 0.521 0.582 ;
      RECT 0.431 0.497 0.481 0.532 ;
      RECT 0.431 0.111 0.481 0.571 ;
    LAYER PO ;
      RECT 0.061 0.071 0.091 1.606 ;
      RECT 0.365 0.069 0.395 1.606 ;
      RECT 0.213 0.071 0.243 1.606 ;
      RECT 1.429 0.065 1.459 1.6 ;
      RECT 1.277 0.065 1.307 1.6 ;
      RECT 0.517 0.071 0.547 1.606 ;
      RECT 0.669 0.069 0.699 1.606 ;
      RECT 1.125 0.069 1.155 1.606 ;
      RECT 0.973 0.069 1.003 1.606 ;
      RECT 0.821 0.069 0.851 1.606 ;
    LAYER NWELL ;
      RECT -0.112 0.679 1.635 1.773 ;
  END
END NBUFFX4_RVT

MACRO AND2X4_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.74 0.553 0.782 ;
      LAYER M1 ;
        RECT 0.553 0.787 0.663 0.815 ;
        RECT 0.491 0.737 0.663 0.787 ;
        RECT 0.553 0.705 0.663 0.737 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.74 0.401 0.782 ;
      LAYER M1 ;
        RECT 0.249 0.787 0.359 0.815 ;
        RECT 0.249 0.737 0.421 0.787 ;
        RECT 0.249 0.705 0.359 0.737 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 ;
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.739 0.15 0.781 0.192 ;
        RECT 1.043 0.15 1.085 0.192 ;
        RECT 1.347 0.152 1.389 0.194 ;
        RECT 0.739 0.242 0.781 0.284 ;
        RECT 1.043 0.242 1.085 0.284 ;
        RECT 1.347 0.244 1.389 0.286 ;
        RECT 0.739 0.334 0.781 0.376 ;
        RECT 1.043 0.334 1.085 0.376 ;
        RECT 1.347 0.336 1.389 0.378 ;
        RECT 0.739 0.426 0.781 0.468 ;
        RECT 1.043 0.426 1.085 0.468 ;
        RECT 1.347 0.428 1.389 0.47 ;
        RECT 0.739 0.838 0.781 0.88 ;
        RECT 1.043 0.838 1.085 0.88 ;
        RECT 1.347 0.838 1.389 0.88 ;
        RECT 0.739 0.93 0.781 0.972 ;
        RECT 1.043 0.93 1.085 0.972 ;
        RECT 1.347 0.93 1.389 0.972 ;
        RECT 0.739 1.022 0.781 1.064 ;
        RECT 1.043 1.022 1.085 1.064 ;
        RECT 1.347 1.022 1.389 1.064 ;
        RECT 0.739 1.114 0.781 1.156 ;
        RECT 1.043 1.114 1.085 1.156 ;
        RECT 1.347 1.114 1.389 1.156 ;
        RECT 0.739 1.206 0.781 1.248 ;
        RECT 1.043 1.206 1.085 1.248 ;
        RECT 1.347 1.206 1.389 1.248 ;
        RECT 0.739 1.298 0.781 1.34 ;
        RECT 1.043 1.298 1.085 1.34 ;
        RECT 1.347 1.298 1.389 1.34 ;
        RECT 0.739 1.39 0.781 1.432 ;
        RECT 1.043 1.39 1.085 1.432 ;
        RECT 1.347 1.39 1.389 1.432 ;
        RECT 0.739 1.482 0.781 1.524 ;
        RECT 1.043 1.482 1.085 1.524 ;
        RECT 1.347 1.482 1.389 1.524 ;
      LAYER M1 ;
        RECT 0.735 0.759 0.785 1.544 ;
        RECT 1.039 0.759 1.089 1.544 ;
        RECT 1.343 0.759 1.393 1.544 ;
        RECT 0.735 0.709 1.478 0.759 ;
        RECT 1.428 0.663 1.478 0.709 ;
        RECT 1.428 0.553 1.575 0.663 ;
        RECT 1.428 0.533 1.478 0.553 ;
        RECT 0.735 0.483 1.478 0.533 ;
        RECT 0.735 0.13 0.785 0.483 ;
        RECT 1.039 0.13 1.089 0.483 ;
        RECT 1.343 0.132 1.393 0.483 ;
    END
    ANTENNADIFFAREA 0.3972 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.891 0.838 0.933 0.88 ;
        RECT 1.195 0.838 1.237 0.88 ;
        RECT 0.891 0.93 0.933 0.972 ;
        RECT 1.195 0.93 1.237 0.972 ;
        RECT 0.891 1.022 0.933 1.064 ;
        RECT 1.195 1.022 1.237 1.064 ;
        RECT 0.891 1.114 0.933 1.156 ;
        RECT 1.195 1.114 1.237 1.156 ;
        RECT 0.891 1.206 0.933 1.248 ;
        RECT 1.195 1.206 1.237 1.248 ;
        RECT 0.435 1.216 0.477 1.258 ;
        RECT 0.891 1.298 0.933 1.34 ;
        RECT 1.195 1.298 1.237 1.34 ;
        RECT 0.435 1.308 0.477 1.35 ;
        RECT 0.891 1.39 0.933 1.432 ;
        RECT 1.195 1.39 1.237 1.432 ;
        RECT 0.435 1.4 0.477 1.442 ;
        RECT 0.891 1.482 0.933 1.524 ;
        RECT 1.195 1.482 1.237 1.524 ;
        RECT 0.435 1.492 0.477 1.534 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.672 1.702 ;
        RECT 0.431 1.196 0.481 1.642 ;
        RECT 0.887 0.818 0.937 1.642 ;
        RECT 1.191 0.818 1.241 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 0.283 0.142 0.325 0.184 ;
        RECT 0.891 0.152 0.933 0.194 ;
        RECT 1.195 0.152 1.237 0.194 ;
        RECT 0.283 0.234 0.325 0.276 ;
        RECT 0.891 0.244 0.933 0.286 ;
        RECT 1.195 0.244 1.237 0.286 ;
        RECT 0.283 0.326 0.325 0.368 ;
        RECT 0.891 0.336 0.933 0.378 ;
        RECT 1.195 0.336 1.237 0.378 ;
        RECT 0.283 0.418 0.325 0.46 ;
      LAYER M1 ;
        RECT 0.279 0.03 0.329 0.48 ;
        RECT 0.887 0.03 0.937 0.398 ;
        RECT 1.191 0.03 1.241 0.398 ;
        RECT 0 -0.03 1.672 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.283 1.308 0.325 1.35 ;
      RECT 0.283 1.216 0.325 1.258 ;
      RECT 0.587 1.308 0.629 1.35 ;
      RECT 0.587 1.4 0.629 1.442 ;
      RECT 0.283 1.492 0.325 1.534 ;
      RECT 0.587 1.492 0.629 1.534 ;
      RECT 0.587 1.216 0.629 1.258 ;
      RECT 0.283 1.4 0.325 1.442 ;
      RECT 1.271 0.595 1.313 0.637 ;
      RECT 0.587 0.234 0.629 0.276 ;
      RECT 0.587 0.418 0.629 0.46 ;
      RECT 0.587 0.326 0.629 0.368 ;
      RECT 0.815 0.595 0.857 0.637 ;
      RECT 1.119 0.595 1.161 0.637 ;
      RECT 0.587 0.142 0.629 0.184 ;
      RECT 0.967 0.595 1.009 0.637 ;
    LAYER M1 ;
      RECT 0.149 0.591 1.333 0.641 ;
      RECT 0.149 0.617 0.199 0.917 ;
      RECT 0.279 0.867 0.329 1.554 ;
      RECT 0.149 0.867 0.633 0.917 ;
      RECT 0.583 0.892 0.633 1.554 ;
      RECT 0.583 0.122 0.633 0.641 ;
    LAYER PO ;
      RECT 0.213 0.071 0.243 1.604 ;
      RECT 0.517 0.071 0.547 1.604 ;
      RECT 0.365 0.071 0.395 1.604 ;
      RECT 0.669 0.071 0.699 1.604 ;
      RECT 0.821 0.072 0.851 1.604 ;
      RECT 1.429 0.072 1.459 1.604 ;
      RECT 1.581 0.072 1.611 1.604 ;
      RECT 1.277 0.072 1.307 1.604 ;
      RECT 1.125 0.072 1.155 1.604 ;
      RECT 0.973 0.072 1.003 1.604 ;
      RECT 0.061 0.071 0.091 1.604 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.787 1.773 ;
  END
END AND2X4_RVT

MACRO NBUFFX8_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.664 0.401 0.706 ;
        RECT 0.511 0.664 0.553 0.706 ;
      LAYER M1 ;
        RECT 0.249 0.71 0.362 0.815 ;
        RECT 0.249 0.66 0.588 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0732 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.739 0.151 0.781 0.193 ;
        RECT 1.043 0.151 1.085 0.193 ;
        RECT 1.347 0.151 1.389 0.193 ;
        RECT 1.651 0.151 1.693 0.193 ;
        RECT 1.955 0.152 1.997 0.194 ;
        RECT 0.739 0.243 0.781 0.285 ;
        RECT 1.043 0.243 1.085 0.285 ;
        RECT 1.347 0.243 1.389 0.285 ;
        RECT 1.651 0.243 1.693 0.285 ;
        RECT 1.955 0.244 1.997 0.286 ;
        RECT 0.739 0.335 0.781 0.377 ;
        RECT 1.043 0.335 1.085 0.377 ;
        RECT 1.347 0.335 1.389 0.377 ;
        RECT 1.651 0.335 1.693 0.377 ;
        RECT 1.955 0.336 1.997 0.378 ;
        RECT 0.739 0.427 0.781 0.469 ;
        RECT 1.043 0.427 1.085 0.469 ;
        RECT 1.347 0.427 1.389 0.469 ;
        RECT 1.651 0.427 1.693 0.469 ;
        RECT 1.955 0.428 1.997 0.47 ;
        RECT 0.739 1.027 0.781 1.069 ;
        RECT 1.043 1.027 1.085 1.069 ;
        RECT 1.347 1.027 1.389 1.069 ;
        RECT 1.651 1.027 1.693 1.069 ;
        RECT 1.955 1.028 1.997 1.07 ;
        RECT 0.739 1.119 0.781 1.161 ;
        RECT 1.043 1.119 1.085 1.161 ;
        RECT 1.347 1.119 1.389 1.161 ;
        RECT 1.651 1.119 1.693 1.161 ;
        RECT 1.955 1.12 1.997 1.162 ;
        RECT 0.739 1.211 0.781 1.253 ;
        RECT 1.043 1.211 1.085 1.253 ;
        RECT 1.347 1.211 1.389 1.253 ;
        RECT 1.651 1.211 1.693 1.253 ;
        RECT 1.955 1.212 1.997 1.254 ;
        RECT 0.739 1.303 0.781 1.345 ;
        RECT 1.043 1.303 1.085 1.345 ;
        RECT 1.347 1.303 1.389 1.345 ;
        RECT 1.651 1.303 1.693 1.345 ;
        RECT 1.955 1.304 1.997 1.346 ;
        RECT 0.739 1.395 0.781 1.437 ;
        RECT 1.043 1.395 1.085 1.437 ;
        RECT 1.347 1.395 1.389 1.437 ;
        RECT 1.651 1.395 1.693 1.437 ;
        RECT 1.955 1.396 1.997 1.438 ;
        RECT 0.739 1.487 0.781 1.529 ;
        RECT 1.043 1.487 1.085 1.529 ;
        RECT 1.347 1.487 1.389 1.529 ;
        RECT 1.651 1.487 1.693 1.529 ;
        RECT 1.955 1.488 1.997 1.53 ;
      LAYER M1 ;
        RECT 1.951 0.942 2.001 1.565 ;
        RECT 0.735 0.942 0.785 1.564 ;
        RECT 1.039 0.942 1.089 1.564 ;
        RECT 1.343 0.942 1.393 1.564 ;
        RECT 1.647 0.942 1.697 1.564 ;
        RECT 0.735 0.892 2.057 0.942 ;
        RECT 2.007 0.663 2.057 0.892 ;
        RECT 2.007 0.587 2.183 0.663 ;
        RECT 0.735 0.537 2.183 0.587 ;
        RECT 0.735 0.116 0.785 0.537 ;
        RECT 1.039 0.116 1.089 0.537 ;
        RECT 1.343 0.116 1.393 0.537 ;
        RECT 1.647 0.116 1.697 0.537 ;
        RECT 1.951 0.117 2.001 0.537 ;
    END
    ANTENNADIFFAREA 0.6952 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.435 1.027 0.477 1.069 ;
        RECT 0.891 1.027 0.933 1.069 ;
        RECT 1.195 1.027 1.237 1.069 ;
        RECT 1.499 1.027 1.541 1.069 ;
        RECT 1.803 1.027 1.845 1.069 ;
        RECT 0.435 1.119 0.477 1.161 ;
        RECT 0.891 1.119 0.933 1.161 ;
        RECT 1.195 1.119 1.237 1.161 ;
        RECT 1.499 1.119 1.541 1.161 ;
        RECT 1.803 1.119 1.845 1.161 ;
        RECT 0.435 1.211 0.477 1.253 ;
        RECT 0.891 1.211 0.933 1.253 ;
        RECT 1.195 1.211 1.237 1.253 ;
        RECT 1.499 1.211 1.541 1.253 ;
        RECT 1.803 1.211 1.845 1.253 ;
        RECT 0.435 1.303 0.477 1.345 ;
        RECT 0.891 1.303 0.933 1.345 ;
        RECT 1.195 1.303 1.237 1.345 ;
        RECT 1.499 1.303 1.541 1.345 ;
        RECT 1.803 1.303 1.845 1.345 ;
        RECT 0.435 1.395 0.477 1.437 ;
        RECT 0.891 1.395 0.933 1.437 ;
        RECT 1.195 1.395 1.237 1.437 ;
        RECT 1.499 1.395 1.541 1.437 ;
        RECT 1.803 1.395 1.845 1.437 ;
        RECT 0.435 1.487 0.477 1.529 ;
        RECT 0.891 1.487 0.933 1.529 ;
        RECT 1.195 1.487 1.237 1.529 ;
        RECT 1.499 1.487 1.541 1.529 ;
        RECT 1.803 1.487 1.845 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 2.28 1.702 ;
        RECT 0.431 0.992 0.481 1.642 ;
        RECT 0.887 0.992 0.937 1.642 ;
        RECT 1.191 0.992 1.241 1.642 ;
        RECT 1.495 0.992 1.545 1.642 ;
        RECT 1.799 0.992 1.849 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 0.435 0.149 0.477 0.191 ;
        RECT 0.891 0.149 0.933 0.191 ;
        RECT 1.195 0.149 1.237 0.191 ;
        RECT 1.499 0.149 1.541 0.191 ;
        RECT 1.803 0.149 1.845 0.191 ;
        RECT 0.435 0.241 0.477 0.283 ;
        RECT 0.891 0.241 0.933 0.283 ;
        RECT 1.195 0.241 1.237 0.283 ;
        RECT 1.499 0.241 1.541 0.283 ;
        RECT 1.803 0.241 1.845 0.283 ;
        RECT 0.435 0.333 0.477 0.375 ;
        RECT 0.891 0.333 0.933 0.375 ;
        RECT 1.195 0.333 1.237 0.375 ;
        RECT 1.499 0.333 1.541 0.375 ;
        RECT 1.803 0.333 1.845 0.375 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.41 ;
        RECT 0.887 0.03 0.937 0.41 ;
        RECT 1.191 0.03 1.241 0.41 ;
        RECT 1.495 0.03 1.545 0.41 ;
        RECT 1.799 0.03 1.849 0.41 ;
        RECT 0 -0.03 2.28 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.283 0.427 0.325 0.469 ;
      RECT 0.283 0.151 0.325 0.193 ;
      RECT 0.815 0.664 0.857 0.706 ;
      RECT 0.967 0.664 1.009 0.706 ;
      RECT 0.283 0.335 0.325 0.377 ;
      RECT 0.283 1.303 0.325 1.345 ;
      RECT 0.283 1.303 0.325 1.345 ;
      RECT 0.283 1.027 0.325 1.069 ;
      RECT 0.283 1.487 0.325 1.529 ;
      RECT 0.587 1.303 0.629 1.345 ;
      RECT 0.283 1.027 0.325 1.069 ;
      RECT 0.283 1.119 0.325 1.161 ;
      RECT 0.283 1.487 0.325 1.529 ;
      RECT 0.283 1.395 0.325 1.437 ;
      RECT 0.283 1.119 0.325 1.161 ;
      RECT 0.283 1.395 0.325 1.437 ;
      RECT 0.587 1.303 0.629 1.345 ;
      RECT 0.587 1.211 0.629 1.253 ;
      RECT 0.587 0.151 0.629 0.193 ;
      RECT 0.587 1.027 0.629 1.069 ;
      RECT 0.587 0.427 0.629 0.469 ;
      RECT 0.587 0.335 0.629 0.377 ;
      RECT 0.587 1.119 0.629 1.161 ;
      RECT 0.587 1.027 0.629 1.069 ;
      RECT 0.587 0.335 0.629 0.377 ;
      RECT 0.587 1.487 0.629 1.529 ;
      RECT 0.587 0.243 0.629 0.285 ;
      RECT 0.587 1.487 0.629 1.529 ;
      RECT 0.587 1.395 0.629 1.437 ;
      RECT 0.587 0.151 0.629 0.193 ;
      RECT 0.587 1.119 0.629 1.161 ;
      RECT 0.587 1.395 0.629 1.437 ;
      RECT 0.587 1.211 0.629 1.253 ;
      RECT 1.879 0.664 1.921 0.706 ;
      RECT 0.283 1.211 0.325 1.253 ;
      RECT 0.283 0.151 0.325 0.193 ;
      RECT 0.283 0.243 0.325 0.285 ;
      RECT 1.575 0.664 1.617 0.706 ;
      RECT 1.727 0.664 1.769 0.706 ;
      RECT 1.423 0.664 1.465 0.706 ;
      RECT 1.271 0.664 1.313 0.706 ;
      RECT 1.119 0.664 1.161 0.706 ;
      RECT 0.283 1.211 0.325 1.253 ;
      RECT 0.283 0.335 0.325 0.377 ;
    LAYER M1 ;
      RECT 0.639 0.66 1.956 0.71 ;
      RECT 0.279 0.892 0.329 1.564 ;
      RECT 0.279 0.502 0.329 0.537 ;
      RECT 0.279 0.116 0.329 0.576 ;
      RECT 0.329 0.939 0.583 0.942 ;
      RECT 0.329 0.931 0.633 0.939 ;
      RECT 0.583 0.892 0.633 1.564 ;
      RECT 0.279 0.892 0.633 0.931 ;
      RECT 0.608 0.892 0.685 0.942 ;
      RECT 0.635 0.85 0.685 0.942 ;
      RECT 0.639 0.609 0.689 0.87 ;
      RECT 0.635 0.537 0.685 0.642 ;
      RECT 0.279 0.537 0.673 0.587 ;
      RECT 0.583 0.116 0.633 0.576 ;
    LAYER PO ;
      RECT 0.061 0.071 0.091 1.606 ;
      RECT 0.517 0.069 0.547 1.606 ;
      RECT 1.885 0.069 1.915 1.606 ;
      RECT 2.037 0.069 2.067 1.606 ;
      RECT 2.189 0.069 2.219 1.606 ;
      RECT 0.213 0.071 0.243 1.606 ;
      RECT 0.365 0.069 0.395 1.606 ;
      RECT 1.733 0.069 1.763 1.606 ;
      RECT 1.581 0.069 1.611 1.606 ;
      RECT 1.429 0.069 1.459 1.606 ;
      RECT 0.669 0.069 0.699 1.606 ;
      RECT 0.821 0.069 0.851 1.606 ;
      RECT 1.277 0.069 1.307 1.606 ;
      RECT 1.125 0.069 1.155 1.606 ;
      RECT 0.973 0.069 1.003 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 2.395 1.773 ;
  END
END NBUFFX8_RVT

MACRO NAND2X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.891 0.553 0.933 ;
      LAYER M1 ;
        RECT 0.553 0.937 0.663 0.967 ;
        RECT 0.456 0.887 0.663 0.937 ;
        RECT 0.553 0.857 0.663 0.887 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.698 0.401 0.74 ;
      LAYER M1 ;
        RECT 0.304 0.664 0.508 0.815 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.195 0.142 1.237 0.184 ;
        RECT 1.195 0.234 1.237 0.276 ;
        RECT 1.195 1.208 1.237 1.25 ;
        RECT 1.195 1.3 1.237 1.342 ;
        RECT 1.195 1.392 1.237 1.434 ;
        RECT 1.195 1.484 1.237 1.526 ;
      LAYER M1 ;
        RECT 1.191 0.969 1.241 1.561 ;
        RECT 1.191 0.861 1.423 0.969 ;
        RECT 1.231 0.857 1.423 0.861 ;
        RECT 1.231 0.505 1.281 0.857 ;
        RECT 1.191 0.455 1.281 0.505 ;
        RECT 1.191 0.114 1.241 0.455 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.739 1.203 0.781 1.245 ;
        RECT 1.043 1.208 1.085 1.25 ;
        RECT 0.435 1.213 0.477 1.255 ;
        RECT 0.739 1.295 0.781 1.337 ;
        RECT 1.043 1.3 1.085 1.342 ;
        RECT 0.435 1.305 0.477 1.347 ;
        RECT 0.739 1.387 0.781 1.429 ;
        RECT 1.043 1.392 1.085 1.434 ;
        RECT 0.435 1.397 0.477 1.439 ;
        RECT 0.739 1.479 0.781 1.521 ;
        RECT 1.043 1.484 1.085 1.526 ;
        RECT 0.435 1.489 0.477 1.531 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.52 1.702 ;
        RECT 0.431 1.193 0.481 1.642 ;
        RECT 0.735 1.183 0.785 1.642 ;
        RECT 1.039 1.188 1.089 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 0.283 0.141 0.325 0.183 ;
        RECT 0.739 0.142 0.781 0.184 ;
        RECT 1.043 0.142 1.085 0.184 ;
        RECT 0.283 0.233 0.325 0.275 ;
        RECT 0.739 0.234 0.781 0.276 ;
        RECT 1.043 0.234 1.085 0.276 ;
        RECT 0.283 0.325 0.325 0.367 ;
        RECT 0.283 0.417 0.325 0.459 ;
      LAYER M1 ;
        RECT 0.279 0.03 0.329 0.479 ;
        RECT 0.735 0.03 0.785 0.296 ;
        RECT 1.039 0.03 1.089 0.296 ;
        RECT 0 -0.03 1.52 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.927 0.642 1.181 0.692 ;
      RECT 0.887 0.906 0.937 1.556 ;
      RECT 0.887 0.455 0.977 0.505 ;
      RECT 0.887 0.114 0.937 0.455 ;
      RECT 0.927 0.692 0.977 0.856 ;
      RECT 0.927 0.505 0.977 0.642 ;
      RECT 0.887 0.856 0.977 0.906 ;
      RECT 0.279 1.07 0.763 1.12 ;
      RECT 0.713 0.781 0.763 1.07 ;
      RECT 0.713 0.731 0.877 0.781 ;
      RECT 0.713 0.663 0.763 0.731 ;
      RECT 0.583 0.613 0.763 0.663 ;
      RECT 0.279 1.12 0.329 1.551 ;
      RECT 0.583 0.106 0.633 0.613 ;
      RECT 0.583 1.12 0.633 1.551 ;
    LAYER PO ;
      RECT 1.125 0.064 1.155 1.607 ;
      RECT 0.821 0.064 0.851 1.602 ;
      RECT 1.429 0.064 1.459 1.6 ;
      RECT 1.277 0.064 1.307 1.605 ;
      RECT 0.973 0.064 1.003 1.6 ;
      RECT 0.061 0.071 0.091 1.601 ;
      RECT 0.213 0.071 0.243 1.601 ;
      RECT 0.517 0.071 0.547 1.601 ;
      RECT 0.365 0.071 0.395 1.601 ;
      RECT 0.669 0.071 0.699 1.601 ;
    LAYER CO ;
      RECT 0.891 1.295 0.933 1.337 ;
      RECT 0.815 0.735 0.857 0.777 ;
      RECT 1.119 0.646 1.161 0.688 ;
      RECT 0.891 0.234 0.933 0.276 ;
      RECT 0.891 0.142 0.933 0.184 ;
      RECT 0.891 0.142 0.933 0.184 ;
      RECT 0.587 0.141 0.629 0.183 ;
      RECT 0.587 0.233 0.629 0.275 ;
      RECT 0.587 0.325 0.629 0.367 ;
      RECT 0.587 0.417 0.629 0.459 ;
      RECT 0.587 1.489 0.629 1.531 ;
      RECT 0.587 1.397 0.629 1.439 ;
      RECT 0.587 1.305 0.629 1.347 ;
      RECT 0.587 1.213 0.629 1.255 ;
      RECT 0.283 1.213 0.325 1.255 ;
      RECT 0.283 1.305 0.325 1.347 ;
      RECT 0.283 1.489 0.325 1.531 ;
      RECT 0.283 1.397 0.325 1.439 ;
      RECT 0.891 1.479 0.933 1.521 ;
      RECT 0.891 1.387 0.933 1.429 ;
      RECT 0.891 1.479 0.933 1.521 ;
      RECT 0.891 1.387 0.933 1.429 ;
      RECT 0.891 1.203 0.933 1.245 ;
      RECT 0.891 1.203 0.933 1.245 ;
      RECT 0.891 1.295 0.933 1.337 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.635 1.781 ;
  END
END NAND2X1_RVT

MACRO NBUFFX2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.216 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.679 0.401 0.721 ;
      LAYER M1 ;
        RECT 0.249 0.725 0.362 0.815 ;
        RECT 0.249 0.675 0.421 0.725 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.587 0.151 0.629 0.193 ;
        RECT 0.891 0.151 0.933 0.193 ;
        RECT 0.587 0.243 0.629 0.285 ;
        RECT 0.891 0.243 0.933 0.285 ;
        RECT 0.587 0.335 0.629 0.377 ;
        RECT 0.891 0.335 0.933 0.377 ;
        RECT 0.587 0.427 0.629 0.469 ;
        RECT 0.891 0.427 0.933 0.469 ;
        RECT 0.587 1.027 0.629 1.069 ;
        RECT 0.891 1.027 0.933 1.069 ;
        RECT 0.587 1.119 0.629 1.161 ;
        RECT 0.891 1.119 0.933 1.161 ;
        RECT 0.587 1.211 0.629 1.253 ;
        RECT 0.891 1.211 0.933 1.253 ;
        RECT 0.587 1.303 0.629 1.345 ;
        RECT 0.891 1.303 0.933 1.345 ;
        RECT 0.587 1.395 0.629 1.437 ;
        RECT 0.891 1.395 0.933 1.437 ;
        RECT 0.587 1.487 0.629 1.529 ;
        RECT 0.891 1.487 0.933 1.529 ;
      LAYER M1 ;
        RECT 0.583 0.942 0.633 1.564 ;
        RECT 0.887 0.942 0.937 1.564 ;
        RECT 0.583 0.892 0.993 0.942 ;
        RECT 0.943 0.663 0.993 0.892 ;
        RECT 0.943 0.587 1.119 0.663 ;
        RECT 0.583 0.537 1.119 0.587 ;
        RECT 0.583 0.116 0.633 0.537 ;
        RECT 0.887 0.116 0.937 0.537 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 0.93 0.325 0.972 ;
        RECT 0.283 1.022 0.325 1.064 ;
        RECT 0.739 1.027 0.781 1.069 ;
        RECT 0.283 1.114 0.325 1.156 ;
        RECT 0.739 1.119 0.781 1.161 ;
        RECT 0.283 1.206 0.325 1.248 ;
        RECT 0.739 1.211 0.781 1.253 ;
        RECT 0.739 1.303 0.781 1.345 ;
        RECT 0.739 1.395 0.781 1.437 ;
        RECT 0.739 1.487 0.781 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.216 1.702 ;
        RECT 0.279 0.91 0.329 1.642 ;
        RECT 0.735 0.992 0.785 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 0.739 0.149 0.781 0.191 ;
        RECT 0.739 0.241 0.781 0.283 ;
        RECT 0.283 0.32 0.325 0.362 ;
        RECT 0.739 0.333 0.781 0.375 ;
        RECT 0.283 0.412 0.325 0.454 ;
        RECT 0.283 0.504 0.325 0.546 ;
      LAYER M1 ;
        RECT 0.279 0.03 0.329 0.567 ;
        RECT 0.735 0.03 0.785 0.41 ;
        RECT 0 -0.03 1.216 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.471 0.66 0.892 0.71 ;
      RECT 0.456 0.887 0.521 0.937 ;
      RECT 0.471 0.532 0.521 0.937 ;
      RECT 0.431 0.887 0.481 1.268 ;
      RECT 0.431 0.887 0.474 0.937 ;
      RECT 0.431 0.3 0.481 0.571 ;
      RECT 0.431 0.532 0.509 0.582 ;
      RECT 0.431 0.497 0.481 0.532 ;
    LAYER PO ;
      RECT 0.061 0.071 0.091 1.606 ;
      RECT 0.365 0.069 0.395 1.606 ;
      RECT 0.213 0.071 0.243 1.606 ;
      RECT 0.517 0.071 0.547 1.606 ;
      RECT 0.669 0.069 0.699 1.606 ;
      RECT 1.125 0.071 1.155 1.606 ;
      RECT 0.973 0.071 1.003 1.606 ;
      RECT 0.821 0.069 0.851 1.606 ;
    LAYER CO ;
      RECT 0.435 1.114 0.477 1.156 ;
      RECT 0.435 1.206 0.477 1.248 ;
      RECT 0.435 0.32 0.477 0.362 ;
      RECT 0.435 0.93 0.477 0.972 ;
      RECT 0.435 1.206 0.477 1.248 ;
      RECT 0.663 0.664 0.705 0.706 ;
      RECT 0.435 1.114 0.477 1.156 ;
      RECT 0.435 1.022 0.477 1.064 ;
      RECT 0.435 0.93 0.477 0.972 ;
      RECT 0.435 0.504 0.477 0.546 ;
      RECT 0.435 0.412 0.477 0.454 ;
      RECT 0.435 0.412 0.477 0.454 ;
      RECT 0.815 0.664 0.857 0.706 ;
      RECT 0.435 1.022 0.477 1.064 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.331 1.773 ;
  END
END NBUFFX2_RVT

MACRO INVX8_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.664 0.401 0.706 ;
        RECT 0.511 0.664 0.553 0.706 ;
        RECT 0.663 0.664 0.705 0.706 ;
        RECT 0.815 0.664 0.857 0.706 ;
        RECT 0.967 0.664 1.009 0.706 ;
        RECT 1.119 0.664 1.161 0.706 ;
        RECT 1.271 0.664 1.313 0.706 ;
        RECT 1.423 0.664 1.465 0.706 ;
      LAYER M1 ;
        RECT 0.249 0.71 0.362 0.815 ;
        RECT 0.249 0.66 1.5 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2928 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.283 0.151 0.325 0.193 ;
        RECT 0.587 0.151 0.629 0.193 ;
        RECT 0.891 0.151 0.933 0.193 ;
        RECT 1.195 0.151 1.237 0.193 ;
        RECT 1.499 0.152 1.541 0.194 ;
        RECT 0.283 0.243 0.325 0.285 ;
        RECT 0.587 0.243 0.629 0.285 ;
        RECT 0.891 0.243 0.933 0.285 ;
        RECT 1.195 0.243 1.237 0.285 ;
        RECT 1.499 0.244 1.541 0.286 ;
        RECT 0.283 0.335 0.325 0.377 ;
        RECT 0.587 0.335 0.629 0.377 ;
        RECT 0.891 0.335 0.933 0.377 ;
        RECT 1.195 0.335 1.237 0.377 ;
        RECT 1.499 0.336 1.541 0.378 ;
        RECT 0.283 0.427 0.325 0.469 ;
        RECT 0.587 0.427 0.629 0.469 ;
        RECT 0.891 0.427 0.933 0.469 ;
        RECT 1.195 0.427 1.237 0.469 ;
        RECT 1.499 0.428 1.541 0.47 ;
        RECT 0.283 1.027 0.325 1.069 ;
        RECT 0.587 1.027 0.629 1.069 ;
        RECT 0.891 1.027 0.933 1.069 ;
        RECT 1.195 1.027 1.237 1.069 ;
        RECT 1.499 1.028 1.541 1.07 ;
        RECT 0.283 1.119 0.325 1.161 ;
        RECT 0.587 1.119 0.629 1.161 ;
        RECT 0.891 1.119 0.933 1.161 ;
        RECT 1.195 1.119 1.237 1.161 ;
        RECT 1.499 1.12 1.541 1.162 ;
        RECT 0.283 1.211 0.325 1.253 ;
        RECT 0.587 1.211 0.629 1.253 ;
        RECT 0.891 1.211 0.933 1.253 ;
        RECT 1.195 1.211 1.237 1.253 ;
        RECT 1.499 1.212 1.541 1.254 ;
        RECT 0.283 1.303 0.325 1.345 ;
        RECT 0.587 1.303 0.629 1.345 ;
        RECT 0.891 1.303 0.933 1.345 ;
        RECT 1.195 1.303 1.237 1.345 ;
        RECT 1.499 1.304 1.541 1.346 ;
        RECT 0.283 1.395 0.325 1.437 ;
        RECT 0.587 1.395 0.629 1.437 ;
        RECT 0.891 1.395 0.933 1.437 ;
        RECT 1.195 1.395 1.237 1.437 ;
        RECT 1.499 1.396 1.541 1.438 ;
        RECT 0.283 1.487 0.325 1.529 ;
        RECT 0.587 1.487 0.629 1.529 ;
        RECT 0.891 1.487 0.933 1.529 ;
        RECT 1.195 1.487 1.237 1.529 ;
        RECT 1.499 1.488 1.541 1.53 ;
      LAYER M1 ;
        RECT 1.495 0.942 1.545 1.565 ;
        RECT 0.279 0.942 0.329 1.564 ;
        RECT 0.583 0.942 0.633 1.564 ;
        RECT 0.887 0.942 0.937 1.564 ;
        RECT 1.191 0.942 1.241 1.564 ;
        RECT 0.279 0.892 1.601 0.942 ;
        RECT 1.551 0.663 1.601 0.892 ;
        RECT 1.551 0.587 1.727 0.663 ;
        RECT 0.279 0.537 1.727 0.587 ;
        RECT 0.279 0.116 0.329 0.537 ;
        RECT 0.583 0.116 0.633 0.537 ;
        RECT 0.887 0.116 0.937 0.537 ;
        RECT 1.191 0.116 1.241 0.537 ;
        RECT 1.495 0.117 1.545 0.537 ;
    END
    ANTENNADIFFAREA 0.6952 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.435 1.027 0.477 1.069 ;
        RECT 0.739 1.027 0.781 1.069 ;
        RECT 1.043 1.027 1.085 1.069 ;
        RECT 1.347 1.027 1.389 1.069 ;
        RECT 0.435 1.119 0.477 1.161 ;
        RECT 0.739 1.119 0.781 1.161 ;
        RECT 1.043 1.119 1.085 1.161 ;
        RECT 1.347 1.119 1.389 1.161 ;
        RECT 0.435 1.211 0.477 1.253 ;
        RECT 0.739 1.211 0.781 1.253 ;
        RECT 1.043 1.211 1.085 1.253 ;
        RECT 1.347 1.211 1.389 1.253 ;
        RECT 0.435 1.303 0.477 1.345 ;
        RECT 0.739 1.303 0.781 1.345 ;
        RECT 1.043 1.303 1.085 1.345 ;
        RECT 1.347 1.303 1.389 1.345 ;
        RECT 0.435 1.395 0.477 1.437 ;
        RECT 0.739 1.395 0.781 1.437 ;
        RECT 1.043 1.395 1.085 1.437 ;
        RECT 1.347 1.395 1.389 1.437 ;
        RECT 0.435 1.487 0.477 1.529 ;
        RECT 0.739 1.487 0.781 1.529 ;
        RECT 1.043 1.487 1.085 1.529 ;
        RECT 1.347 1.487 1.389 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.824 1.702 ;
        RECT 0.431 0.992 0.481 1.642 ;
        RECT 0.735 0.992 0.785 1.642 ;
        RECT 1.039 0.992 1.089 1.642 ;
        RECT 1.343 0.992 1.393 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 0.435 0.149 0.477 0.191 ;
        RECT 0.739 0.149 0.781 0.191 ;
        RECT 1.043 0.149 1.085 0.191 ;
        RECT 1.347 0.149 1.389 0.191 ;
        RECT 0.435 0.241 0.477 0.283 ;
        RECT 0.739 0.241 0.781 0.283 ;
        RECT 1.043 0.241 1.085 0.283 ;
        RECT 1.347 0.241 1.389 0.283 ;
        RECT 0.435 0.333 0.477 0.375 ;
        RECT 0.739 0.333 0.781 0.375 ;
        RECT 1.043 0.333 1.085 0.375 ;
        RECT 1.347 0.333 1.389 0.375 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.41 ;
        RECT 0.735 0.03 0.785 0.41 ;
        RECT 1.039 0.03 1.089 0.41 ;
        RECT 1.343 0.03 1.393 0.41 ;
        RECT 0 -0.03 1.824 0.03 ;
    END
  END VSS
  OBS
    LAYER PO ;
      RECT 1.429 0.069 1.459 1.606 ;
      RECT 1.581 0.069 1.611 1.606 ;
      RECT 1.733 0.069 1.763 1.606 ;
      RECT 1.277 0.069 1.307 1.606 ;
      RECT 1.125 0.069 1.155 1.606 ;
      RECT 0.973 0.069 1.003 1.606 ;
      RECT 0.213 0.069 0.243 1.606 ;
      RECT 0.365 0.069 0.395 1.606 ;
      RECT 0.821 0.069 0.851 1.606 ;
      RECT 0.669 0.069 0.699 1.606 ;
      RECT 0.517 0.069 0.547 1.606 ;
      RECT 0.061 0.069 0.091 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.939 1.773 ;
  END
END INVX8_RVT

MACRO AOI221X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.879 0.401 0.921 ;
      LAYER M1 ;
        RECT 0.249 0.857 0.404 0.967 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.601 0.553 0.643 ;
      LAYER M1 ;
        RECT 0.401 0.553 0.555 0.663 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.136 0.857 0.178 ;
      LAYER M1 ;
        RECT 0.705 0.097 0.863 0.207 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.875 0.705 0.917 ;
      LAYER M1 ;
        RECT 0.553 1.009 0.663 1.119 ;
        RECT 0.613 0.921 0.663 1.009 ;
        RECT 0.613 0.871 0.725 0.921 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.119 0.777 1.161 0.819 ;
      LAYER M1 ;
        RECT 1.007 0.773 1.181 0.823 ;
        RECT 1.009 0.705 1.119 0.773 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0201 ;
  END A5
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.803 0.134 1.845 0.176 ;
        RECT 1.803 0.226 1.845 0.268 ;
        RECT 1.803 0.318 1.845 0.36 ;
        RECT 1.803 0.411 1.845 0.453 ;
        RECT 1.803 0.858 1.845 0.9 ;
        RECT 1.803 0.95 1.845 0.992 ;
        RECT 1.803 1.042 1.845 1.084 ;
        RECT 1.803 1.134 1.845 1.176 ;
        RECT 1.803 1.226 1.845 1.268 ;
        RECT 1.803 1.318 1.845 1.36 ;
        RECT 1.803 1.41 1.845 1.452 ;
      LAYER M1 ;
        RECT 1.799 1.271 1.849 1.472 ;
        RECT 1.769 1.161 1.879 1.271 ;
        RECT 1.799 0.853 1.849 1.161 ;
        RECT 1.799 0.852 1.889 0.853 ;
        RECT 1.799 0.803 1.899 0.852 ;
        RECT 1.849 0.476 1.899 0.803 ;
        RECT 1.799 0.426 1.899 0.476 ;
        RECT 1.799 0.114 1.849 0.426 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.347 1.225 1.389 1.267 ;
        RECT 1.651 1.226 1.693 1.268 ;
        RECT 1.347 1.317 1.389 1.359 ;
        RECT 1.651 1.318 1.693 1.36 ;
        RECT 0.435 1.407 0.477 1.449 ;
        RECT 1.347 1.409 1.389 1.451 ;
        RECT 1.651 1.41 1.693 1.452 ;
        RECT 0.435 1.499 0.477 1.541 ;
        RECT 1.347 1.501 1.389 1.543 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 2.128 1.702 ;
        RECT 0.431 1.387 0.481 1.642 ;
        RECT 1.343 1.167 1.393 1.642 ;
        RECT 1.647 1.206 1.697 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 1.651 0.134 1.693 0.176 ;
        RECT 1.651 0.226 1.693 0.268 ;
        RECT 0.587 0.265 0.629 0.307 ;
        RECT 1.043 0.272 1.085 0.314 ;
        RECT 1.651 0.318 1.693 0.36 ;
        RECT 1.347 0.335 1.389 0.377 ;
        RECT 0.587 0.357 0.629 0.399 ;
        RECT 1.651 0.411 1.693 0.453 ;
        RECT 1.347 0.427 1.389 0.469 ;
      LAYER M1 ;
        RECT 1.343 0.03 1.393 0.489 ;
        RECT 1.647 0.03 1.697 0.473 ;
        RECT 0.583 0.03 0.633 0.419 ;
        RECT 1.04 0.03 1.09 0.334 ;
        RECT 0 -0.03 2.128 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.283 1.509 0.325 1.551 ;
      RECT 0.739 1.175 0.781 1.217 ;
      RECT 0.739 1.083 0.781 1.125 ;
      RECT 0.587 1.509 0.629 1.551 ;
      RECT 0.587 1.325 0.629 1.367 ;
      RECT 0.283 0.353 0.325 0.395 ;
      RECT 1.043 1.233 1.085 1.275 ;
      RECT 0.891 0.374 0.933 0.416 ;
      RECT 0.891 1.509 0.933 1.551 ;
      RECT 1.043 1.141 1.085 1.183 ;
      RECT 0.891 0.282 0.933 0.324 ;
      RECT 0.283 0.261 0.325 0.303 ;
      RECT 0.891 1.325 0.933 1.367 ;
      RECT 1.195 1.509 1.237 1.551 ;
      RECT 1.195 1.325 1.237 1.367 ;
      RECT 1.043 1.509 1.085 1.551 ;
      RECT 1.195 1.141 1.237 1.183 ;
      RECT 1.195 0.28 1.237 0.322 ;
      RECT 1.043 1.325 1.085 1.367 ;
      RECT 1.043 1.417 1.085 1.459 ;
      RECT 0.587 1.417 0.629 1.459 ;
      RECT 0.891 1.417 0.933 1.459 ;
      RECT 1.499 0.335 1.541 0.377 ;
      RECT 1.727 0.627 1.769 0.669 ;
      RECT 1.423 0.8 1.465 0.842 ;
      RECT 1.499 0.427 1.541 0.469 ;
      RECT 1.195 1.417 1.237 1.459 ;
      RECT 1.499 1.409 1.541 1.451 ;
      RECT 1.499 1.501 1.541 1.543 ;
      RECT 1.499 1.317 1.541 1.359 ;
      RECT 1.499 1.225 1.541 1.267 ;
      RECT 1.195 1.233 1.237 1.275 ;
      RECT 0.283 1.325 0.325 1.367 ;
      RECT 0.283 1.417 0.325 1.459 ;
    LAYER M1 ;
      RECT 1.419 0.774 1.469 0.907 ;
      RECT 0.887 0.908 1.469 0.957 ;
      RECT 1.233 0.907 1.469 0.908 ;
      RECT 0.279 0.241 0.329 0.731 ;
      RECT 0.887 0.781 0.937 0.908 ;
      RECT 0.279 0.731 0.937 0.781 ;
      RECT 0.887 0.262 0.937 0.731 ;
      RECT 1.191 0.253 1.241 0.673 ;
      RECT 1.191 0.673 1.282 0.674 ;
      RECT 1.191 0.674 1.283 0.723 ;
      RECT 1.191 1.081 1.241 1.571 ;
      RECT 1.191 1.031 1.283 1.081 ;
      RECT 1.233 0.958 1.283 1.031 ;
      RECT 0.887 0.957 1.283 0.958 ;
      RECT 1.233 0.723 1.283 0.907 ;
      RECT 1.495 0.623 1.789 0.673 ;
      RECT 1.495 1.002 1.665 1.052 ;
      RECT 1.615 0.673 1.665 1.002 ;
      RECT 1.495 1.052 1.545 1.563 ;
      RECT 1.495 1.001 1.545 1.002 ;
      RECT 1.495 0.315 1.545 0.623 ;
      RECT 0.735 1.021 1.089 1.071 ;
      RECT 1.039 1.071 1.089 1.571 ;
      RECT 0.735 1.071 0.785 1.237 ;
      RECT 0.583 1.337 0.633 1.571 ;
      RECT 0.279 1.287 0.937 1.337 ;
      RECT 0.887 1.337 0.937 1.571 ;
      RECT 0.279 1.337 0.329 1.571 ;
    LAYER PO ;
      RECT 1.885 0.063 1.915 1.604 ;
      RECT 1.581 0.063 1.611 1.604 ;
      RECT 1.277 0.075 1.307 1.621 ;
      RECT 1.733 0.064 1.763 1.604 ;
      RECT 1.429 0.059 1.459 1.621 ;
      RECT 2.037 0.063 2.067 1.604 ;
      RECT 0.669 0.072 0.699 1.621 ;
      RECT 0.517 0.072 0.547 1.621 ;
      RECT 0.365 0.067 0.395 1.621 ;
      RECT 0.061 0.072 0.091 1.621 ;
      RECT 0.973 0.076 1.003 1.621 ;
      RECT 0.821 0.072 0.851 1.621 ;
      RECT 0.213 0.072 0.243 1.621 ;
      RECT 1.125 0.076 1.155 1.621 ;
    LAYER NWELL ;
      RECT -0.115 0.679 2.243 1.773 ;
  END
END AOI221X1_RVT

MACRO INVX4_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.216 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.664 0.401 0.706 ;
        RECT 0.511 0.664 0.553 0.706 ;
        RECT 0.663 0.664 0.705 0.706 ;
        RECT 0.815 0.664 0.857 0.706 ;
      LAYER M1 ;
        RECT 0.249 0.71 0.362 0.815 ;
        RECT 0.249 0.66 0.892 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1464 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.283 0.151 0.325 0.193 ;
        RECT 0.587 0.151 0.629 0.193 ;
        RECT 0.891 0.151 0.933 0.193 ;
        RECT 0.283 0.243 0.325 0.285 ;
        RECT 0.587 0.243 0.629 0.285 ;
        RECT 0.891 0.243 0.933 0.285 ;
        RECT 0.283 0.335 0.325 0.377 ;
        RECT 0.587 0.335 0.629 0.377 ;
        RECT 0.891 0.335 0.933 0.377 ;
        RECT 0.283 0.427 0.325 0.469 ;
        RECT 0.587 0.427 0.629 0.469 ;
        RECT 0.891 0.427 0.933 0.469 ;
        RECT 0.283 1.027 0.325 1.069 ;
        RECT 0.587 1.027 0.629 1.069 ;
        RECT 0.891 1.027 0.933 1.069 ;
        RECT 0.283 1.119 0.325 1.161 ;
        RECT 0.587 1.119 0.629 1.161 ;
        RECT 0.891 1.119 0.933 1.161 ;
        RECT 0.283 1.211 0.325 1.253 ;
        RECT 0.587 1.211 0.629 1.253 ;
        RECT 0.891 1.211 0.933 1.253 ;
        RECT 0.283 1.303 0.325 1.345 ;
        RECT 0.587 1.303 0.629 1.345 ;
        RECT 0.891 1.303 0.933 1.345 ;
        RECT 0.283 1.395 0.325 1.437 ;
        RECT 0.587 1.395 0.629 1.437 ;
        RECT 0.891 1.395 0.933 1.437 ;
        RECT 0.283 1.487 0.325 1.529 ;
        RECT 0.587 1.487 0.629 1.529 ;
        RECT 0.891 1.487 0.933 1.529 ;
      LAYER M1 ;
        RECT 0.279 0.942 0.329 1.564 ;
        RECT 0.583 0.942 0.633 1.564 ;
        RECT 0.887 0.942 0.937 1.564 ;
        RECT 0.279 0.892 0.992 0.942 ;
        RECT 0.942 0.663 0.992 0.892 ;
        RECT 0.942 0.587 1.119 0.663 ;
        RECT 0.279 0.537 1.119 0.587 ;
        RECT 0.279 0.116 0.329 0.537 ;
        RECT 0.583 0.116 0.633 0.537 ;
        RECT 0.887 0.116 0.937 0.537 ;
    END
    ANTENNADIFFAREA 0.3976 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.435 1.027 0.477 1.069 ;
        RECT 0.739 1.027 0.781 1.069 ;
        RECT 0.435 1.119 0.477 1.161 ;
        RECT 0.739 1.119 0.781 1.161 ;
        RECT 0.435 1.211 0.477 1.253 ;
        RECT 0.739 1.211 0.781 1.253 ;
        RECT 0.435 1.303 0.477 1.345 ;
        RECT 0.739 1.303 0.781 1.345 ;
        RECT 0.435 1.395 0.477 1.437 ;
        RECT 0.739 1.395 0.781 1.437 ;
        RECT 0.435 1.487 0.477 1.529 ;
        RECT 0.739 1.487 0.781 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.216 1.702 ;
        RECT 0.431 0.992 0.481 1.642 ;
        RECT 0.735 0.992 0.785 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 0.435 0.149 0.477 0.191 ;
        RECT 0.739 0.149 0.781 0.191 ;
        RECT 0.435 0.241 0.477 0.283 ;
        RECT 0.739 0.241 0.781 0.283 ;
        RECT 0.435 0.333 0.477 0.375 ;
        RECT 0.739 0.333 0.781 0.375 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.41 ;
        RECT 0.735 0.03 0.785 0.41 ;
        RECT 0 -0.03 1.216 0.03 ;
    END
  END VSS
  OBS
    LAYER PO ;
      RECT 1.125 0.065 1.155 1.6 ;
      RECT 0.973 0.065 1.003 1.6 ;
      RECT 0.213 0.071 0.243 1.606 ;
      RECT 0.365 0.069 0.395 1.606 ;
      RECT 0.821 0.069 0.851 1.606 ;
      RECT 0.669 0.069 0.699 1.606 ;
      RECT 0.517 0.069 0.547 1.606 ;
      RECT 0.061 0.071 0.091 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.331 1.773 ;
  END
END INVX4_RVT

MACRO XNOR2X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.967 0.61 1.009 0.652 ;
        RECT 1.879 0.675 1.921 0.717 ;
      LAYER M1 ;
        RECT 0.962 0.672 1.941 0.722 ;
        RECT 0.962 0.553 1.119 0.672 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0405 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.745 0.705 0.787 ;
        RECT 1.575 0.807 1.617 0.849 ;
      LAYER M1 ;
        RECT 0.658 0.803 1.655 0.853 ;
        RECT 0.658 0.705 0.815 0.803 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0378 ;
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 2.259 0.183 2.301 0.225 ;
        RECT 2.259 0.275 2.301 0.317 ;
        RECT 2.259 0.367 2.301 0.409 ;
        RECT 2.259 0.459 2.301 0.501 ;
        RECT 2.259 0.961 2.301 1.003 ;
        RECT 2.259 1.073 2.301 1.115 ;
        RECT 2.259 1.165 2.301 1.207 ;
        RECT 2.259 1.257 2.301 1.299 ;
        RECT 2.259 1.349 2.301 1.391 ;
        RECT 2.259 1.441 2.301 1.483 ;
      LAYER M1 ;
        RECT 2.255 0.967 2.305 1.546 ;
        RECT 2.255 0.917 2.487 0.967 ;
        RECT 2.31 0.857 2.487 0.917 ;
        RECT 2.31 0.554 2.36 0.857 ;
        RECT 2.255 0.504 2.36 0.554 ;
        RECT 2.255 0.148 2.305 0.504 ;
    END
    ANTENNADIFFAREA 0.1234 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 2.107 0.849 2.149 0.891 ;
        RECT 2.107 0.941 2.149 0.983 ;
        RECT 2.107 1.033 2.149 1.075 ;
        RECT 2.107 1.125 2.149 1.167 ;
        RECT 0.283 1.149 0.325 1.191 ;
        RECT 2.107 1.217 2.149 1.259 ;
        RECT 0.283 1.241 0.325 1.283 ;
        RECT 0.587 1.253 0.629 1.295 ;
        RECT 1.043 1.253 1.085 1.295 ;
        RECT 1.651 1.253 1.693 1.295 ;
        RECT 2.107 1.309 2.149 1.351 ;
        RECT 0.283 1.333 0.325 1.375 ;
        RECT 2.107 1.401 2.149 1.443 ;
        RECT 2.107 1.493 2.149 1.535 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 2.584 1.702 ;
        RECT 0.279 1.129 0.329 1.642 ;
        RECT 0.583 1.218 0.633 1.642 ;
        RECT 1.039 1.218 1.089 1.642 ;
        RECT 1.647 1.218 1.697 1.642 ;
        RECT 2.103 0.814 2.153 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.107 0.17 2.149 0.212 ;
        RECT 2.107 0.262 2.149 0.304 ;
        RECT 0.587 0.274 0.629 0.316 ;
        RECT 1.043 0.274 1.085 0.316 ;
        RECT 1.651 0.274 1.693 0.316 ;
        RECT 0.283 0.275 0.325 0.317 ;
        RECT 2.107 0.354 2.149 0.396 ;
        RECT 2.107 0.446 2.149 0.488 ;
      LAYER M1 ;
        RECT 0.279 0.371 0.612 0.421 ;
        RECT 0.562 0.32 0.612 0.371 ;
        RECT 0.562 0.27 1.12 0.32 ;
        RECT 1.616 0.27 1.785 0.32 ;
        RECT 2.103 0.03 2.153 0.526 ;
        RECT 0.279 0.03 0.329 0.371 ;
        RECT 1.735 0.03 1.785 0.27 ;
        RECT 0 -0.03 2.584 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 1.499 1.243 1.541 1.285 ;
      RECT 1.955 0.367 1.997 0.409 ;
      RECT 1.955 1.073 1.997 1.115 ;
      RECT 2.183 0.608 2.225 0.65 ;
      RECT 1.347 1.012 1.389 1.054 ;
      RECT 1.955 0.275 1.997 0.317 ;
      RECT 0.435 1.243 0.477 1.285 ;
      RECT 1.955 0.367 1.997 0.409 ;
      RECT 1.803 1.243 1.845 1.285 ;
      RECT 0.891 0.985 0.933 1.027 ;
      RECT 0.739 1.022 0.781 1.064 ;
      RECT 1.195 1.243 1.237 1.285 ;
      RECT 1.955 0.961 1.997 1.003 ;
      RECT 0.359 0.608 0.401 0.65 ;
      RECT 1.955 0.961 1.997 1.003 ;
      RECT 1.955 1.073 1.997 1.115 ;
      RECT 1.803 0.375 1.845 0.417 ;
      RECT 0.739 0.39 0.781 0.432 ;
      RECT 1.347 0.329 1.389 0.371 ;
      RECT 1.955 1.174 1.997 1.216 ;
      RECT 0.435 0.275 0.477 0.317 ;
      RECT 0.891 0.412 0.933 0.454 ;
      RECT 1.271 0.576 1.313 0.618 ;
      RECT 1.499 0.375 1.541 0.417 ;
      RECT 1.195 0.264 1.237 0.306 ;
    LAYER M1 ;
      RECT 0.355 1.018 0.816 1.068 ;
      RECT 0.735 0.37 0.785 0.471 ;
      RECT 0.355 0.471 0.785 0.521 ;
      RECT 0.324 0.604 0.405 0.654 ;
      RECT 0.355 0.521 0.405 0.604 ;
      RECT 0.355 0.654 0.405 1.018 ;
      RECT 0.846 0.408 1.224 0.458 ;
      RECT 1.174 0.458 1.224 0.572 ;
      RECT 1.174 0.572 1.35 0.622 ;
      RECT 0.48 0.571 0.896 0.621 ;
      RECT 0.48 0.918 0.937 0.968 ;
      RECT 0.887 0.968 0.937 1.068 ;
      RECT 0.846 0.458 0.896 0.571 ;
      RECT 0.48 0.621 0.53 0.918 ;
      RECT 1.991 0.604 2.26 0.654 ;
      RECT 1.36 0.375 1.41 0.471 ;
      RECT 1.327 0.325 1.41 0.375 ;
      RECT 1.951 0.24 2.001 0.471 ;
      RECT 1.991 0.654 2.041 0.809 ;
      RECT 1.951 0.809 2.041 0.859 ;
      RECT 1.951 1.058 2.001 1.305 ;
      RECT 1.312 1.008 2.001 1.058 ;
      RECT 1.951 0.859 2.001 1.008 ;
      RECT 1.991 0.521 2.041 0.604 ;
      RECT 1.36 0.471 2.041 0.521 ;
      RECT 0.462 0.153 1.241 0.203 ;
      RECT 1.191 0.203 1.241 0.326 ;
      RECT 0.4 0.271 0.512 0.321 ;
      RECT 0.462 0.203 0.512 0.271 ;
      RECT 1.464 0.371 1.88 0.421 ;
      RECT 1.16 1.239 1.576 1.289 ;
      RECT 0.431 1.118 1.849 1.168 ;
      RECT 1.799 1.168 1.849 1.32 ;
      RECT 0.431 1.168 0.481 1.32 ;
    LAYER PO ;
      RECT 0.365 0.066 0.395 1.606 ;
      RECT 1.581 0.066 1.611 1.606 ;
      RECT 0.517 0.066 0.547 1.606 ;
      RECT 1.429 0.068 1.459 1.606 ;
      RECT 2.493 0.068 2.523 1.606 ;
      RECT 0.061 0.068 0.091 1.606 ;
      RECT 0.669 0.068 0.699 1.606 ;
      RECT 0.213 0.068 0.243 1.606 ;
      RECT 0.821 0.068 0.851 1.606 ;
      RECT 1.733 0.068 1.763 1.606 ;
      RECT 1.125 0.068 1.155 1.606 ;
      RECT 2.037 0.068 2.067 1.606 ;
      RECT 0.973 0.068 1.003 1.606 ;
      RECT 2.189 0.068 2.219 1.606 ;
      RECT 2.341 0.068 2.371 1.606 ;
      RECT 1.277 0.068 1.307 1.606 ;
      RECT 1.885 0.068 1.915 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 2.699 1.781 ;
  END
END XNOR2X1_RVT

MACRO OR4X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.666 0.401 0.708 ;
      LAYER M1 ;
        RECT 0.249 0.662 0.421 0.712 ;
        RECT 0.249 0.553 0.359 0.662 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.666 0.553 0.708 ;
      LAYER M1 ;
        RECT 0.507 0.857 0.663 0.967 ;
        RECT 0.507 0.646 0.557 0.857 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.666 0.705 0.708 ;
      LAYER M1 ;
        RECT 0.659 0.511 0.709 0.728 ;
        RECT 0.659 0.401 0.815 0.511 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.666 0.857 0.708 ;
      LAYER M1 ;
        RECT 0.811 0.705 0.967 0.815 ;
        RECT 0.811 0.646 0.861 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A4
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.803 0.148 1.845 0.19 ;
        RECT 1.803 0.242 1.845 0.284 ;
        RECT 1.803 0.334 1.845 0.376 ;
        RECT 1.803 0.427 1.845 0.469 ;
        RECT 1.803 0.823 1.845 0.865 ;
        RECT 1.803 0.915 1.845 0.957 ;
        RECT 1.803 1.009 1.845 1.051 ;
        RECT 1.803 1.101 1.845 1.143 ;
        RECT 1.803 1.194 1.845 1.236 ;
        RECT 1.803 1.286 1.845 1.328 ;
        RECT 1.803 1.38 1.845 1.422 ;
        RECT 1.803 1.472 1.845 1.514 ;
      LAYER M1 ;
        RECT 1.799 0.812 1.849 1.549 ;
        RECT 1.799 0.762 1.969 0.812 ;
        RECT 1.919 0.489 1.969 0.762 ;
        RECT 1.799 0.439 1.969 0.489 ;
        RECT 1.799 0.128 1.849 0.439 ;
        RECT 1.919 0.359 1.969 0.439 ;
        RECT 1.919 0.249 2.031 0.359 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 0.833 0.325 0.875 ;
        RECT 0.283 0.93 0.325 0.972 ;
        RECT 1.347 0.931 1.389 0.973 ;
        RECT 0.283 1.024 0.325 1.066 ;
        RECT 1.347 1.024 1.389 1.066 ;
        RECT 1.043 1.085 1.085 1.127 ;
        RECT 0.283 1.116 0.325 1.158 ;
        RECT 1.347 1.116 1.389 1.158 ;
        RECT 1.651 1.116 1.693 1.158 ;
        RECT 0.283 1.209 0.325 1.251 ;
        RECT 1.347 1.209 1.389 1.251 ;
        RECT 1.651 1.209 1.693 1.251 ;
        RECT 0.283 1.301 0.325 1.343 ;
        RECT 1.347 1.301 1.389 1.343 ;
        RECT 1.651 1.301 1.693 1.343 ;
        RECT 0.283 1.395 0.325 1.437 ;
        RECT 1.347 1.395 1.389 1.437 ;
        RECT 1.651 1.395 1.693 1.437 ;
        RECT 0.283 1.487 0.325 1.529 ;
        RECT 1.347 1.487 1.389 1.529 ;
        RECT 1.651 1.487 1.693 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 2.128 1.702 ;
        RECT 0.279 0.813 0.329 1.642 ;
        RECT 1.039 1.065 1.089 1.642 ;
        RECT 1.343 0.911 1.393 1.642 ;
        RECT 1.647 1.096 1.697 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 1.043 0.141 1.085 0.183 ;
        RECT 1.347 0.141 1.389 0.183 ;
        RECT 1.651 0.141 1.693 0.183 ;
        RECT 0.435 0.179 0.477 0.221 ;
        RECT 0.739 0.179 0.781 0.221 ;
        RECT 1.347 0.233 1.389 0.275 ;
        RECT 1.651 0.233 1.693 0.275 ;
        RECT 1.347 0.325 1.389 0.367 ;
        RECT 1.651 0.325 1.693 0.367 ;
      LAYER M1 ;
        RECT 1.343 0.03 1.393 0.387 ;
        RECT 1.647 0.03 1.697 0.387 ;
        RECT 0.431 0.03 0.481 0.241 ;
        RECT 0.735 0.03 0.785 0.241 ;
        RECT 1.039 0.03 1.089 0.203 ;
        RECT 0 -0.03 2.128 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 1.499 0.334 1.541 0.376 ;
      RECT 1.499 0.242 1.541 0.284 ;
      RECT 1.499 0.148 1.541 0.19 ;
      RECT 1.499 0.427 1.541 0.469 ;
      RECT 1.499 1.458 1.541 1.5 ;
      RECT 1.499 1.366 1.541 1.408 ;
      RECT 1.423 0.667 1.465 0.709 ;
      RECT 1.499 1.272 1.541 1.314 ;
      RECT 1.499 1.18 1.541 1.222 ;
      RECT 1.499 1.087 1.541 1.129 ;
      RECT 1.499 0.995 1.541 1.037 ;
      RECT 1.499 0.901 1.541 0.943 ;
      RECT 0.891 0.23 0.933 0.272 ;
      RECT 0.283 0.23 0.325 0.272 ;
      RECT 0.891 1.473 0.933 1.515 ;
      RECT 0.891 1.381 0.933 1.423 ;
      RECT 0.891 1.287 0.933 1.329 ;
      RECT 0.891 1.195 0.933 1.237 ;
      RECT 0.891 1.102 0.933 1.144 ;
      RECT 0.587 0.23 0.629 0.272 ;
      RECT 0.891 1.01 0.933 1.052 ;
      RECT 1.195 0.812 1.237 0.854 ;
      RECT 0.891 0.918 0.933 0.96 ;
      RECT 1.119 0.67 1.161 0.712 ;
      RECT 1.195 0.245 1.237 0.287 ;
      RECT 1.195 0.151 1.237 0.193 ;
      RECT 1.195 1.09 1.237 1.132 ;
      RECT 1.195 0.998 1.237 1.04 ;
      RECT 1.195 0.904 1.237 0.946 ;
      RECT 1.727 0.667 1.769 0.709 ;
    LAYER M1 ;
      RECT 1.029 0.666 1.181 0.716 ;
      RECT 1.029 0.341 1.079 0.666 ;
      RECT 0.279 0.291 1.079 0.341 ;
      RECT 1.029 0.716 1.079 0.898 ;
      RECT 0.887 0.898 1.079 0.948 ;
      RECT 0.887 0.209 0.937 0.291 ;
      RECT 0.887 0.948 0.937 1.55 ;
      RECT 0.279 0.21 0.329 0.291 ;
      RECT 0.583 0.21 0.633 0.291 ;
      RECT 1.34 0.663 1.485 0.713 ;
      RECT 1.34 0.552 1.39 0.663 ;
      RECT 1.192 0.527 1.39 0.552 ;
      RECT 1.191 0.502 1.39 0.527 ;
      RECT 1.34 0.713 1.39 0.803 ;
      RECT 1.191 0.803 1.39 0.853 ;
      RECT 1.191 0.853 1.241 1.152 ;
      RECT 1.191 0.792 1.241 0.803 ;
      RECT 1.191 0.131 1.241 0.502 ;
      RECT 1.495 0.897 1.665 0.947 ;
      RECT 1.615 0.663 1.789 0.713 ;
      RECT 1.615 0.552 1.665 0.663 ;
      RECT 1.495 0.502 1.665 0.552 ;
      RECT 1.615 0.713 1.665 0.897 ;
      RECT 1.495 0.947 1.545 1.535 ;
      RECT 1.495 0.881 1.545 0.897 ;
      RECT 1.495 0.128 1.545 0.502 ;
    LAYER PO ;
      RECT 1.125 0.071 1.155 1.612 ;
      RECT 1.277 0.071 1.307 1.612 ;
      RECT 1.429 0.071 1.459 1.61 ;
      RECT 1.581 0.072 1.611 1.61 ;
      RECT 0.973 0.072 1.003 1.61 ;
      RECT 0.061 0.072 0.091 1.61 ;
      RECT 2.037 0.072 2.067 1.61 ;
      RECT 0.821 0.072 0.851 1.61 ;
      RECT 1.885 0.072 1.915 1.61 ;
      RECT 1.733 0.071 1.763 1.61 ;
      RECT 0.213 0.072 0.243 1.61 ;
      RECT 0.669 0.072 0.699 1.61 ;
      RECT 0.365 0.072 0.395 1.61 ;
      RECT 0.517 0.072 0.547 1.61 ;
    LAYER NWELL ;
      RECT -0.115 0.679 2.243 1.801 ;
  END
END OR4X1_RVT

MACRO INVX1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.664 0.401 0.706 ;
      LAYER M1 ;
        RECT 0.249 0.71 0.362 0.815 ;
        RECT 0.249 0.66 0.421 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.283 0.151 0.325 0.193 ;
        RECT 0.283 0.243 0.325 0.285 ;
        RECT 0.283 0.335 0.325 0.377 ;
        RECT 0.283 0.427 0.325 0.469 ;
        RECT 0.283 1.027 0.325 1.069 ;
        RECT 0.283 1.119 0.325 1.161 ;
        RECT 0.283 1.211 0.325 1.253 ;
        RECT 0.283 1.303 0.325 1.345 ;
        RECT 0.283 1.395 0.325 1.437 ;
        RECT 0.283 1.487 0.325 1.529 ;
      LAYER M1 ;
        RECT 0.279 0.942 0.329 1.564 ;
        RECT 0.279 0.892 0.521 0.942 ;
        RECT 0.471 0.663 0.521 0.892 ;
        RECT 0.471 0.587 0.663 0.663 ;
        RECT 0.279 0.537 0.663 0.587 ;
        RECT 0.279 0.116 0.329 0.537 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.435 1.027 0.477 1.069 ;
        RECT 0.435 1.119 0.477 1.161 ;
        RECT 0.435 1.211 0.477 1.253 ;
        RECT 0.435 1.303 0.477 1.345 ;
        RECT 0.435 1.395 0.477 1.437 ;
        RECT 0.435 1.487 0.477 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 0.76 1.702 ;
        RECT 0.431 0.992 0.481 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.435 0.149 0.477 0.191 ;
        RECT 0.435 0.241 0.477 0.283 ;
        RECT 0.435 0.333 0.477 0.375 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.41 ;
        RECT 0 -0.03 0.76 0.03 ;
    END
  END VSS
  OBS
    LAYER PO ;
      RECT 0.213 0.071 0.243 1.606 ;
      RECT 0.365 0.069 0.395 1.606 ;
      RECT 0.669 0.071 0.699 1.606 ;
      RECT 0.517 0.071 0.547 1.606 ;
      RECT 0.061 0.071 0.091 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 0.875 1.773 ;
  END
END INVX1_RVT

MACRO OR3X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.667 0.401 0.709 ;
      LAYER M1 ;
        RECT 0.249 0.705 0.405 0.815 ;
        RECT 0.355 0.647 0.405 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.667 0.553 0.709 ;
      LAYER M1 ;
        RECT 0.507 0.857 0.663 0.967 ;
        RECT 0.507 0.647 0.557 0.857 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.667 0.705 0.709 ;
      LAYER M1 ;
        RECT 0.66 0.553 0.815 0.729 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END A3
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.043 0.151 1.085 0.193 ;
        RECT 1.043 0.245 1.085 0.287 ;
        RECT 1.043 0.337 1.085 0.379 ;
        RECT 1.043 0.43 1.085 0.472 ;
        RECT 1.043 0.823 1.085 0.865 ;
        RECT 1.043 0.915 1.085 0.957 ;
        RECT 1.043 1.009 1.085 1.051 ;
        RECT 1.043 1.101 1.085 1.143 ;
        RECT 1.043 1.194 1.085 1.236 ;
        RECT 1.043 1.286 1.085 1.328 ;
        RECT 1.043 1.38 1.085 1.422 ;
        RECT 1.043 1.472 1.085 1.514 ;
      LAYER M1 ;
        RECT 1.039 0.853 1.089 1.534 ;
        RECT 1.039 0.803 1.244 0.853 ;
        RECT 1.194 0.476 1.244 0.803 ;
        RECT 1.039 0.476 1.089 0.492 ;
        RECT 1.039 0.426 1.244 0.476 ;
        RECT 1.039 0.131 1.089 0.426 ;
        RECT 1.194 0.359 1.244 0.426 ;
        RECT 1.161 0.249 1.271 0.359 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 0.931 0.325 0.973 ;
        RECT 0.891 0.932 0.933 0.974 ;
        RECT 0.283 1.024 0.325 1.066 ;
        RECT 0.891 1.024 0.933 1.066 ;
        RECT 0.283 1.116 0.325 1.158 ;
        RECT 0.891 1.116 0.933 1.158 ;
        RECT 0.283 1.209 0.325 1.251 ;
        RECT 0.891 1.209 0.933 1.251 ;
        RECT 0.283 1.301 0.325 1.343 ;
        RECT 0.891 1.301 0.933 1.343 ;
        RECT 0.283 1.395 0.325 1.437 ;
        RECT 0.891 1.395 0.933 1.437 ;
        RECT 0.283 1.487 0.325 1.529 ;
        RECT 0.891 1.487 0.933 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.52 1.702 ;
        RECT 0.279 0.911 0.329 1.642 ;
        RECT 0.887 0.912 0.937 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 0.891 0.141 0.933 0.183 ;
        RECT 0.891 0.233 0.933 0.275 ;
        RECT 0.435 0.262 0.477 0.304 ;
        RECT 0.739 0.262 0.781 0.304 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.324 ;
        RECT 0.735 0.03 0.785 0.324 ;
        RECT 0.887 0.03 0.937 0.295 ;
        RECT 0 -0.03 1.52 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.279 0.374 0.931 0.424 ;
      RECT 0.881 0.399 0.931 0.852 ;
      RECT 0.735 0.802 0.906 0.852 ;
      RECT 0.901 0.663 1.029 0.713 ;
      RECT 0.735 0.818 0.785 1.549 ;
      RECT 0.279 0.317 0.329 0.399 ;
      RECT 0.583 0.317 0.633 0.399 ;
    LAYER PO ;
      RECT 0.973 0.071 1.003 1.609 ;
      RECT 1.125 0.071 1.155 1.609 ;
      RECT 1.277 0.071 1.307 1.609 ;
      RECT 0.061 0.071 0.091 1.609 ;
      RECT 0.821 0.071 0.851 1.609 ;
      RECT 0.213 0.071 0.243 1.609 ;
      RECT 0.669 0.071 0.699 1.609 ;
      RECT 0.365 0.071 0.395 1.609 ;
      RECT 0.517 0.071 0.547 1.609 ;
    LAYER CO ;
      RECT 0.967 0.667 1.009 0.709 ;
      RECT 0.739 0.838 0.781 0.88 ;
      RECT 0.283 0.337 0.325 0.379 ;
      RECT 0.739 1.487 0.781 1.529 ;
      RECT 0.739 1.395 0.781 1.437 ;
      RECT 0.739 1.301 0.781 1.343 ;
      RECT 0.739 1.209 0.781 1.251 ;
      RECT 0.739 1.116 0.781 1.158 ;
      RECT 0.587 0.337 0.629 0.379 ;
      RECT 0.739 1.024 0.781 1.066 ;
      RECT 0.739 0.93 0.781 0.972 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.635 1.773 ;
  END
END OR3X1_RVT

MACRO OR2X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.216 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.662 0.401 0.704 ;
      LAYER M1 ;
        RECT 0.249 0.857 0.405 0.967 ;
        RECT 0.355 0.642 0.405 0.857 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0303 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.662 0.553 0.704 ;
      LAYER M1 ;
        RECT 0.502 0.642 0.663 0.815 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0303 ;
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.891 0.219 0.933 0.261 ;
        RECT 0.891 0.311 0.933 0.353 ;
        RECT 0.891 0.403 0.933 0.445 ;
        RECT 0.891 0.495 0.933 0.537 ;
        RECT 0.891 0.836 0.933 0.878 ;
        RECT 0.891 0.928 0.933 0.97 ;
        RECT 0.891 1.02 0.933 1.062 ;
        RECT 0.891 1.112 0.933 1.154 ;
        RECT 0.891 1.204 0.933 1.246 ;
        RECT 0.891 1.296 0.933 1.338 ;
        RECT 0.891 1.39 0.933 1.432 ;
        RECT 0.891 1.482 0.933 1.524 ;
      LAYER M1 ;
        RECT 0.887 0.866 0.937 1.544 ;
        RECT 0.887 0.816 1.043 0.866 ;
        RECT 0.993 0.558 1.043 0.816 ;
        RECT 0.887 0.511 1.043 0.558 ;
        RECT 0.887 0.508 1.119 0.511 ;
        RECT 0.887 0.199 0.937 0.508 ;
        RECT 0.993 0.401 1.119 0.508 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.107 0.325 1.149 ;
        RECT 0.739 1.107 0.781 1.149 ;
        RECT 0.283 1.2 0.325 1.242 ;
        RECT 0.739 1.2 0.781 1.242 ;
        RECT 0.283 1.292 0.325 1.334 ;
        RECT 0.739 1.292 0.781 1.334 ;
        RECT 0.283 1.386 0.325 1.428 ;
        RECT 0.739 1.386 0.781 1.428 ;
        RECT 0.283 1.478 0.325 1.52 ;
        RECT 0.739 1.478 0.781 1.52 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.216 1.702 ;
        RECT 0.279 1.087 0.329 1.642 ;
        RECT 0.735 1.086 0.785 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 0.739 0.147 0.781 0.189 ;
        RECT 0.739 0.239 0.781 0.281 ;
        RECT 0.739 0.331 0.781 0.373 ;
        RECT 0.435 0.334 0.477 0.376 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.399 ;
        RECT 0.735 0.03 0.785 0.393 ;
        RECT 0 -0.03 1.216 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.742 0.658 0.889 0.708 ;
      RECT 0.726 0.486 0.776 0.956 ;
      RECT 0.279 0.297 0.329 0.512 ;
      RECT 0.582 0.905 0.732 0.955 ;
      RECT 0.583 0.889 0.633 1.525 ;
      RECT 0.278 0.486 0.733 0.536 ;
      RECT 0.583 0.299 0.633 0.512 ;
    LAYER PO ;
      RECT 1.125 0.073 1.155 1.6 ;
      RECT 0.973 0.073 1.003 1.6 ;
      RECT 0.061 0.073 0.091 1.604 ;
      RECT 0.821 0.073 0.851 1.604 ;
      RECT 0.213 0.073 0.243 1.604 ;
      RECT 0.669 0.073 0.699 1.604 ;
      RECT 0.365 0.073 0.395 1.604 ;
      RECT 0.517 0.073 0.547 1.604 ;
    LAYER CO ;
      RECT 0.815 0.662 0.857 0.704 ;
      RECT 0.587 0.909 0.629 0.951 ;
      RECT 0.587 1.001 0.629 1.043 ;
      RECT 0.283 0.409 0.325 0.451 ;
      RECT 0.283 0.317 0.325 0.359 ;
      RECT 0.587 1.463 0.629 1.505 ;
      RECT 0.587 1.371 0.629 1.413 ;
      RECT 0.587 1.277 0.629 1.319 ;
      RECT 0.587 1.185 0.629 1.227 ;
      RECT 0.587 0.319 0.629 0.361 ;
      RECT 0.587 1.093 0.629 1.135 ;
      RECT 0.587 0.411 0.629 0.453 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.331 1.773 ;
  END
END OR2X1_RVT

MACRO MUX21X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.615 0.401 0.657 ;
      LAYER M1 ;
        RECT 0.355 0.663 0.405 0.692 ;
        RECT 0.249 0.553 0.415 0.663 ;
        RECT 0.355 0.499 0.405 0.553 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0189 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.271 1.042 1.313 1.084 ;
      LAYER M1 ;
        RECT 1.251 1.009 1.423 1.119 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0189 ;
  END A2
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.119 0.634 1.161 0.676 ;
        RECT 0.815 0.733 0.857 0.775 ;
        RECT 0.511 1.077 0.553 1.119 ;
      LAYER M1 ;
        RECT 0.507 0.779 0.557 1.154 ;
        RECT 0.811 0.779 0.967 0.815 ;
        RECT 0.507 0.729 0.967 0.779 ;
        RECT 0.811 0.705 0.967 0.729 ;
        RECT 0.917 0.664 0.967 0.705 ;
        RECT 1.115 0.664 1.165 0.696 ;
        RECT 0.917 0.614 1.165 0.664 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0378 ;
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.651 0.187 1.693 0.229 ;
        RECT 1.651 0.279 1.693 0.321 ;
        RECT 1.651 0.371 1.693 0.413 ;
        RECT 1.651 0.463 1.693 0.505 ;
        RECT 1.651 0.873 1.693 0.915 ;
        RECT 1.651 0.965 1.693 1.007 ;
        RECT 1.651 1.077 1.693 1.119 ;
        RECT 1.651 1.169 1.693 1.211 ;
        RECT 1.651 1.261 1.693 1.303 ;
        RECT 1.651 1.353 1.693 1.395 ;
        RECT 1.651 1.445 1.693 1.487 ;
      LAYER M1 ;
        RECT 1.647 0.815 1.697 1.55 ;
        RECT 1.647 0.765 1.88 0.815 ;
        RECT 1.751 0.705 1.88 0.765 ;
        RECT 1.751 0.558 1.801 0.705 ;
        RECT 1.647 0.508 1.801 0.558 ;
        RECT 1.647 0.152 1.697 0.508 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.587 1.405 0.629 1.447 ;
        RECT 0.891 1.405 0.933 1.447 ;
        RECT 1.043 1.405 1.085 1.447 ;
        RECT 1.499 1.405 1.541 1.447 ;
        RECT 0.587 1.497 0.629 1.539 ;
        RECT 0.891 1.497 0.933 1.539 ;
        RECT 1.043 1.497 1.085 1.539 ;
        RECT 1.499 1.497 1.541 1.539 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.976 1.702 ;
        RECT 0.583 1.385 0.633 1.642 ;
        RECT 0.887 1.385 0.937 1.642 ;
        RECT 1.039 1.385 1.089 1.642 ;
        RECT 1.495 1.385 1.545 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 0.587 0.141 0.629 0.183 ;
        RECT 0.891 0.142 0.933 0.184 ;
        RECT 1.043 0.142 1.085 0.184 ;
        RECT 1.499 0.174 1.541 0.216 ;
        RECT 0.587 0.233 0.629 0.275 ;
        RECT 0.891 0.234 0.933 0.276 ;
        RECT 1.043 0.234 1.085 0.276 ;
        RECT 1.499 0.266 1.541 0.308 ;
        RECT 1.499 0.358 1.541 0.4 ;
        RECT 1.499 0.45 1.541 0.492 ;
      LAYER M1 ;
        RECT 1.495 0.03 1.545 0.558 ;
        RECT 0.887 0.03 0.937 0.296 ;
        RECT 1.039 0.03 1.089 0.296 ;
        RECT 0.583 0.03 0.633 0.295 ;
        RECT 0 -0.03 1.976 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.283 1.38 0.325 1.422 ;
      RECT 1.347 0.266 1.389 0.308 ;
      RECT 0.283 1.472 0.325 1.514 ;
      RECT 0.283 1.38 0.325 1.422 ;
      RECT 1.119 1.047 1.161 1.089 ;
      RECT 1.347 0.174 1.389 0.216 ;
      RECT 0.283 0.265 0.325 0.307 ;
      RECT 1.347 1.481 1.389 1.523 ;
      RECT 0.283 0.173 0.325 0.215 ;
      RECT 1.575 0.612 1.617 0.654 ;
      RECT 0.739 1.17 0.781 1.212 ;
      RECT 0.739 0.181 0.781 0.223 ;
      RECT 0.283 1.196 0.325 1.238 ;
      RECT 1.347 1.389 1.389 1.431 ;
      RECT 1.347 1.389 1.389 1.431 ;
      RECT 0.739 0.273 0.781 0.315 ;
      RECT 1.347 1.481 1.389 1.523 ;
      RECT 0.283 1.288 0.325 1.33 ;
      RECT 0.283 1.288 0.325 1.33 ;
      RECT 0.511 0.451 0.553 0.493 ;
      RECT 0.283 1.472 0.325 1.514 ;
    LAYER M1 ;
      RECT 1.115 0.752 1.293 0.802 ;
      RECT 0.507 0.514 1.293 0.564 ;
      RECT 1.243 0.564 1.293 0.752 ;
      RECT 0.735 1.074 1.165 1.124 ;
      RECT 1.115 0.802 1.165 1.074 ;
      RECT 0.507 0.424 0.557 0.514 ;
      RECT 0.735 1.124 0.785 1.232 ;
      RECT 0.735 0.161 0.785 0.514 ;
      RECT 1.343 0.608 1.652 0.658 ;
      RECT 0.279 1.285 1.564 1.335 ;
      RECT 1.514 0.658 1.564 1.285 ;
      RECT 0.149 0.337 0.199 0.894 ;
      RECT 0.149 0.287 0.329 0.337 ;
      RECT 0.279 0.138 0.329 0.287 ;
      RECT 0.279 1.335 0.329 1.549 ;
      RECT 0.279 0.944 0.329 1.285 ;
      RECT 0.149 0.894 0.329 0.944 ;
      RECT 1.343 1.335 1.393 1.55 ;
      RECT 1.343 0.139 1.393 0.608 ;
    LAYER PO ;
      RECT 1.125 0.072 1.155 0.711 ;
      RECT 0.061 0.071 0.091 1.609 ;
      RECT 0.365 0.069 0.395 1.609 ;
      RECT 0.213 0.071 0.243 1.609 ;
      RECT 1.581 0.072 1.611 1.61 ;
      RECT 1.733 0.072 1.763 1.61 ;
      RECT 1.885 0.072 1.915 1.61 ;
      RECT 0.669 0.071 0.699 1.609 ;
      RECT 0.517 0.071 0.547 0.525 ;
      RECT 0.821 0.072 0.851 1.61 ;
      RECT 1.125 1.015 1.155 1.61 ;
      RECT 0.973 0.072 1.003 1.61 ;
      RECT 1.277 0.072 1.307 1.61 ;
      RECT 1.429 0.072 1.459 1.61 ;
      RECT 0.517 1.045 0.547 1.609 ;
    LAYER NWELL ;
      RECT -0.115 0.679 2.091 1.773 ;
  END
END MUX21X1_RVT

MACRO OAI22X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.271 0.81 0.421 0.817 ;
        RECT 0.249 0.71 0.421 0.81 ;
        RECT 0.249 0.701 0.359 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0276 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.482 0.553 1.524 ;
      LAYER M1 ;
        RECT 0.401 1.571 0.511 1.576 ;
        RECT 0.401 1.461 0.573 1.571 ;
        RECT 0.426 1.46 0.573 1.461 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0276 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.744 0.857 0.786 ;
      LAYER M1 ;
        RECT 0.811 1.002 0.968 1.139 ;
        RECT 0.811 0.715 0.861 1.002 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0276 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.747 0.705 0.789 ;
      LAYER M1 ;
        RECT 0.56 0.963 0.709 0.986 ;
        RECT 0.553 0.854 0.709 0.963 ;
        RECT 0.659 0.723 0.709 0.854 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0276 ;
  END A4
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.499 0.239 1.541 0.281 ;
        RECT 1.499 0.331 1.541 0.373 ;
        RECT 1.499 0.423 1.541 0.465 ;
        RECT 1.499 0.987 1.541 1.029 ;
        RECT 1.499 1.079 1.541 1.121 ;
        RECT 1.499 1.171 1.541 1.213 ;
        RECT 1.499 1.263 1.541 1.305 ;
        RECT 1.499 1.355 1.541 1.397 ;
      LAYER M1 ;
        RECT 1.495 1.006 1.545 1.426 ;
        RECT 1.495 0.956 1.684 1.006 ;
        RECT 1.634 0.542 1.684 0.956 ;
        RECT 1.495 0.53 1.684 0.542 ;
        RECT 1.495 0.492 1.759 0.53 ;
        RECT 1.495 0.188 1.545 0.492 ;
        RECT 1.599 0.392 1.759 0.492 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.079 0.325 1.121 ;
        RECT 0.283 1.171 0.325 1.213 ;
        RECT 1.347 1.171 1.389 1.213 ;
        RECT 0.283 1.263 0.325 1.305 ;
        RECT 1.347 1.263 1.389 1.305 ;
        RECT 0.283 1.355 0.325 1.397 ;
        RECT 0.891 1.355 0.933 1.397 ;
        RECT 1.347 1.355 1.389 1.397 ;
        RECT 1.043 1.392 1.085 1.434 ;
        RECT 1.043 1.484 1.085 1.526 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.824 1.702 ;
        RECT 0.279 0.958 0.329 1.642 ;
        RECT 0.887 1.335 0.937 1.642 ;
        RECT 1.039 1.363 1.089 1.642 ;
        RECT 1.343 1.133 1.393 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.043 0.143 1.085 0.185 ;
        RECT 1.347 0.203 1.389 0.245 ;
        RECT 1.043 0.235 1.085 0.277 ;
        RECT 0.435 0.239 0.477 0.281 ;
        RECT 1.347 0.295 1.389 0.337 ;
        RECT 1.043 0.327 1.085 0.369 ;
        RECT 0.435 0.331 0.477 0.373 ;
        RECT 0.435 0.423 0.477 0.465 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.512 ;
        RECT 1.039 0.03 1.089 0.404 ;
        RECT 1.343 0.03 1.393 0.399 ;
        RECT 0 -0.03 1.824 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.383 0.681 1.469 0.699 ;
      RECT 1.383 0.613 1.469 0.631 ;
      RECT 1.231 0.631 1.469 0.681 ;
      RECT 1.231 0.681 1.281 0.956 ;
      RECT 1.231 0.542 1.281 0.631 ;
      RECT 1.191 1.006 1.241 1.426 ;
      RECT 1.191 0.956 1.281 1.006 ;
      RECT 1.191 0.188 1.241 0.492 ;
      RECT 1.191 0.492 1.281 0.542 ;
      RECT 1.079 0.664 1.165 0.75 ;
      RECT 1.079 0.75 1.129 1.226 ;
      RECT 0.583 1.226 1.129 1.276 ;
      RECT 1.079 0.616 1.129 0.664 ;
      RECT 0.735 0.566 1.129 0.616 ;
      RECT 0.735 0.212 0.785 0.566 ;
      RECT 0.583 1.276 0.633 1.393 ;
      RECT 0.583 1.106 0.633 1.226 ;
      RECT 0.583 0.095 0.937 0.145 ;
      RECT 0.279 0.598 0.633 0.648 ;
      RECT 0.583 0.145 0.633 0.598 ;
      RECT 0.887 0.145 0.937 0.504 ;
      RECT 0.279 0.178 0.329 0.598 ;
    LAYER PO ;
      RECT 0.061 0.101 0.091 1.469 ;
      RECT 0.517 0.101 0.547 1.567 ;
      RECT 0.213 0.101 0.243 1.469 ;
      RECT 0.973 0.101 1.003 1.469 ;
      RECT 0.821 0.101 0.851 1.469 ;
      RECT 0.669 0.101 0.699 1.469 ;
      RECT 1.125 0.054 1.155 1.608 ;
      RECT 1.429 0.069 1.459 1.608 ;
      RECT 1.277 0.101 1.307 1.469 ;
      RECT 0.365 0.101 0.395 1.469 ;
      RECT 1.581 0.101 1.611 1.469 ;
      RECT 1.733 0.101 1.763 1.469 ;
    LAYER CO ;
      RECT 0.587 1.23 0.629 1.272 ;
      RECT 0.587 1.138 0.629 1.18 ;
      RECT 0.587 1.322 0.629 1.364 ;
      RECT 0.587 0.423 0.629 0.465 ;
      RECT 1.195 0.239 1.237 0.281 ;
      RECT 0.891 0.331 0.933 0.373 ;
      RECT 0.891 0.239 0.933 0.281 ;
      RECT 1.195 0.331 1.237 0.373 ;
      RECT 0.739 0.331 0.781 0.373 ;
      RECT 1.119 0.686 1.161 0.728 ;
      RECT 0.283 0.423 0.325 0.465 ;
      RECT 0.283 0.331 0.325 0.373 ;
      RECT 0.891 0.423 0.933 0.465 ;
      RECT 0.739 0.239 0.781 0.281 ;
      RECT 0.739 0.423 0.781 0.465 ;
      RECT 0.283 0.239 0.325 0.281 ;
      RECT 0.587 0.331 0.629 0.373 ;
      RECT 1.195 1.079 1.237 1.121 ;
      RECT 1.195 1.171 1.237 1.213 ;
      RECT 1.195 1.263 1.237 1.305 ;
      RECT 1.195 1.355 1.237 1.397 ;
      RECT 0.587 0.239 0.629 0.281 ;
      RECT 1.423 0.635 1.465 0.677 ;
    LAYER NWELL ;
      RECT -0.135 0.679 1.94 1.787 ;
  END
END OAI22X1_RVT

MACRO NOR4X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.665 0.401 0.707 ;
      LAYER M1 ;
        RECT 0.355 0.663 0.405 0.747 ;
        RECT 0.249 0.553 0.405 0.663 ;
        RECT 0.355 0.551 0.405 0.553 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.665 0.553 0.707 ;
      LAYER M1 ;
        RECT 0.401 0.95 0.511 0.967 ;
        RECT 0.401 0.857 0.557 0.95 ;
        RECT 0.507 0.645 0.557 0.857 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.665 0.705 0.707 ;
      LAYER M1 ;
        RECT 0.553 1.009 0.719 1.119 ;
        RECT 0.659 0.645 0.709 1.009 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.665 0.857 0.707 ;
      LAYER M1 ;
        RECT 0.809 0.645 0.967 0.815 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A4
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.499 0.148 1.541 0.19 ;
        RECT 1.499 0.242 1.541 0.284 ;
        RECT 1.499 0.334 1.541 0.376 ;
        RECT 1.499 0.427 1.541 0.469 ;
        RECT 1.499 0.912 1.541 0.954 ;
        RECT 1.499 1.006 1.541 1.048 ;
        RECT 1.499 1.098 1.541 1.14 ;
        RECT 1.499 1.191 1.541 1.233 ;
        RECT 1.499 1.283 1.541 1.325 ;
        RECT 1.499 1.377 1.541 1.419 ;
        RECT 1.499 1.469 1.541 1.511 ;
      LAYER M1 ;
        RECT 1.495 0.942 1.545 1.531 ;
        RECT 1.495 0.892 1.699 0.942 ;
        RECT 1.649 0.511 1.699 0.892 ;
        RECT 1.617 0.487 1.727 0.511 ;
        RECT 1.495 0.487 1.545 0.489 ;
        RECT 1.495 0.437 1.727 0.487 ;
        RECT 1.495 0.128 1.545 0.437 ;
        RECT 1.617 0.401 1.727 0.437 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 0.93 0.325 0.972 ;
        RECT 1.043 0.997 1.085 1.039 ;
        RECT 0.283 1.024 0.325 1.066 ;
        RECT 1.043 1.089 1.085 1.131 ;
        RECT 1.347 1.113 1.389 1.155 ;
        RECT 0.283 1.116 0.325 1.158 ;
        RECT 1.043 1.181 1.085 1.223 ;
        RECT 1.347 1.206 1.389 1.248 ;
        RECT 0.283 1.209 0.325 1.251 ;
        RECT 1.347 1.298 1.389 1.34 ;
        RECT 0.283 1.301 0.325 1.343 ;
        RECT 1.347 1.392 1.389 1.434 ;
        RECT 0.283 1.395 0.325 1.437 ;
        RECT 1.347 1.484 1.389 1.526 ;
        RECT 0.283 1.487 0.325 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.824 1.702 ;
        RECT 0.279 0.91 0.329 1.642 ;
        RECT 1.039 0.977 1.089 1.642 ;
        RECT 1.343 1.093 1.393 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.347 0.148 1.389 0.19 ;
        RECT 1.043 0.149 1.085 0.191 ;
        RECT 1.043 0.241 1.085 0.283 ;
        RECT 1.347 0.242 1.389 0.284 ;
        RECT 0.435 0.269 0.477 0.311 ;
        RECT 0.739 0.28 0.781 0.322 ;
        RECT 1.347 0.334 1.389 0.376 ;
      LAYER M1 ;
        RECT 1.343 0.03 1.393 0.396 ;
        RECT 0.735 0.03 0.785 0.342 ;
        RECT 0.431 0.03 0.481 0.331 ;
        RECT 1.039 0.03 1.089 0.303 ;
        RECT 0 -0.03 1.824 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.279 0.397 1.083 0.447 ;
      RECT 0.887 0.872 1.083 0.922 ;
      RECT 1.033 0.747 1.181 0.797 ;
      RECT 1.033 0.447 1.083 0.747 ;
      RECT 1.033 0.797 1.083 0.872 ;
      RECT 0.279 0.261 0.329 0.397 ;
      RECT 0.583 0.261 0.633 0.397 ;
      RECT 0.887 0.26 0.937 0.397 ;
      RECT 0.887 0.922 0.937 1.535 ;
      RECT 1.191 0.498 1.365 0.548 ;
      RECT 1.192 0.851 1.365 0.876 ;
      RECT 1.191 0.876 1.365 0.901 ;
      RECT 1.314 0.661 1.485 0.711 ;
      RECT 1.314 0.548 1.364 0.661 ;
      RECT 1.314 0.711 1.364 0.851 ;
      RECT 1.191 0.128 1.241 0.498 ;
      RECT 1.191 0.901 1.241 1.224 ;
    LAYER PO ;
      RECT 1.429 0.068 1.459 1.609 ;
      RECT 1.581 0.068 1.611 1.609 ;
      RECT 1.125 0.068 1.155 1.609 ;
      RECT 1.277 0.068 1.307 1.609 ;
      RECT 0.973 0.068 1.003 1.609 ;
      RECT 1.733 0.072 1.763 1.609 ;
      RECT 0.061 0.072 0.091 1.609 ;
      RECT 0.821 0.072 0.851 1.609 ;
      RECT 0.213 0.072 0.243 1.609 ;
      RECT 0.669 0.072 0.699 1.609 ;
      RECT 0.365 0.072 0.395 1.609 ;
      RECT 0.517 0.072 0.547 1.609 ;
    LAYER CO ;
      RECT 0.891 1.458 0.933 1.5 ;
      RECT 0.891 1.366 0.933 1.408 ;
      RECT 0.891 1.272 0.933 1.314 ;
      RECT 0.891 1.18 0.933 1.222 ;
      RECT 1.423 0.665 1.465 0.707 ;
      RECT 1.195 1.07 1.237 1.112 ;
      RECT 1.195 0.978 1.237 1.02 ;
      RECT 0.891 1.087 0.933 1.129 ;
      RECT 0.587 0.281 0.629 0.323 ;
      RECT 0.891 0.995 0.933 1.037 ;
      RECT 1.195 0.884 1.237 0.926 ;
      RECT 1.195 1.162 1.237 1.204 ;
      RECT 1.119 0.751 1.161 0.793 ;
      RECT 1.195 0.242 1.237 0.284 ;
      RECT 1.195 0.148 1.237 0.19 ;
      RECT 0.891 0.28 0.933 0.322 ;
      RECT 0.283 0.281 0.325 0.323 ;
      RECT 0.891 0.903 0.933 0.945 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.939 1.773 ;
  END
END NOR4X1_RVT

MACRO NOR2X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.665 0.401 0.707 ;
      LAYER M1 ;
        RECT 0.249 0.631 0.421 0.815 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0303 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.665 0.553 0.707 ;
      LAYER M1 ;
        RECT 0.489 0.553 0.663 0.733 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0303 ;
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.195 0.151 1.237 0.193 ;
        RECT 1.195 0.245 1.237 0.287 ;
        RECT 1.195 0.337 1.237 0.379 ;
        RECT 1.195 0.43 1.237 0.472 ;
        RECT 1.195 0.841 1.237 0.883 ;
        RECT 1.195 0.933 1.237 0.975 ;
        RECT 1.195 1.027 1.237 1.069 ;
        RECT 1.195 1.119 1.237 1.161 ;
        RECT 1.195 1.212 1.237 1.254 ;
        RECT 1.195 1.304 1.237 1.346 ;
        RECT 1.195 1.398 1.237 1.44 ;
        RECT 1.195 1.49 1.237 1.532 ;
      LAYER M1 ;
        RECT 1.191 0.824 1.241 1.552 ;
        RECT 1.191 0.774 1.395 0.824 ;
        RECT 1.345 0.511 1.395 0.774 ;
        RECT 1.313 0.49 1.423 0.511 ;
        RECT 1.191 0.49 1.241 0.492 ;
        RECT 1.191 0.44 1.423 0.49 ;
        RECT 1.191 0.131 1.241 0.44 ;
        RECT 1.313 0.401 1.423 0.44 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 0.931 0.325 0.973 ;
        RECT 1.043 0.931 1.085 0.973 ;
        RECT 0.739 1.008 0.781 1.05 ;
        RECT 0.283 1.024 0.325 1.066 ;
        RECT 1.043 1.024 1.085 1.066 ;
        RECT 0.739 1.1 0.781 1.142 ;
        RECT 0.283 1.116 0.325 1.158 ;
        RECT 1.043 1.116 1.085 1.158 ;
        RECT 0.283 1.209 0.325 1.251 ;
        RECT 1.043 1.209 1.085 1.251 ;
        RECT 0.283 1.301 0.325 1.343 ;
        RECT 1.043 1.301 1.085 1.343 ;
        RECT 0.283 1.395 0.325 1.437 ;
        RECT 1.043 1.395 1.085 1.437 ;
        RECT 0.283 1.487 0.325 1.529 ;
        RECT 1.043 1.487 1.085 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.52 1.702 ;
        RECT 0.279 0.911 0.329 1.642 ;
        RECT 0.735 0.988 0.785 1.642 ;
        RECT 1.039 0.911 1.089 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 0.739 0.141 0.781 0.183 ;
        RECT 1.043 0.141 1.085 0.183 ;
        RECT 0.435 0.176 0.477 0.218 ;
        RECT 0.739 0.233 0.781 0.275 ;
        RECT 1.043 0.233 1.085 0.275 ;
        RECT 0.435 0.268 0.477 0.31 ;
        RECT 1.043 0.325 1.085 0.367 ;
      LAYER M1 ;
        RECT 1.039 0.03 1.089 0.387 ;
        RECT 0.431 0.03 0.481 0.33 ;
        RECT 0.735 0.03 0.785 0.295 ;
        RECT 0 -0.03 1.52 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.279 0.383 0.775 0.433 ;
      RECT 0.583 0.813 0.775 0.863 ;
      RECT 0.725 0.666 0.877 0.716 ;
      RECT 0.725 0.433 0.775 0.666 ;
      RECT 0.725 0.716 0.775 0.813 ;
      RECT 0.279 0.174 0.329 0.383 ;
      RECT 0.583 0.174 0.633 0.383 ;
      RECT 0.583 0.863 0.633 1.552 ;
      RECT 0.887 0.773 1.06 0.823 ;
      RECT 0.887 0.502 1.061 0.552 ;
      RECT 1.01 0.711 1.06 0.773 ;
      RECT 1.01 0.661 1.181 0.711 ;
      RECT 1.01 0.552 1.06 0.661 ;
      RECT 0.887 0.823 0.937 1.152 ;
      RECT 0.887 0.131 0.937 0.502 ;
    LAYER PO ;
      RECT 1.125 0.071 1.155 1.612 ;
      RECT 1.277 0.071 1.307 1.612 ;
      RECT 0.821 0.071 0.851 1.612 ;
      RECT 0.973 0.071 1.003 1.612 ;
      RECT 0.061 0.071 0.091 1.612 ;
      RECT 1.429 0.071 1.459 1.612 ;
      RECT 0.213 0.071 0.243 1.612 ;
      RECT 0.669 0.071 0.699 1.612 ;
      RECT 0.365 0.071 0.395 1.612 ;
      RECT 0.517 0.071 0.547 1.612 ;
    LAYER CO ;
      RECT 0.587 1.49 0.629 1.532 ;
      RECT 0.587 1.396 0.629 1.438 ;
      RECT 0.587 1.304 0.629 1.346 ;
      RECT 0.587 1.211 0.629 1.253 ;
      RECT 0.587 0.194 0.629 0.236 ;
      RECT 0.283 0.194 0.325 0.236 ;
      RECT 0.891 0.812 0.933 0.854 ;
      RECT 0.587 0.842 0.629 0.884 ;
      RECT 0.587 0.934 0.629 0.976 ;
      RECT 0.587 1.027 0.629 1.069 ;
      RECT 0.815 0.67 0.857 0.712 ;
      RECT 0.891 0.245 0.933 0.287 ;
      RECT 0.891 0.151 0.933 0.193 ;
      RECT 1.119 0.665 1.161 0.707 ;
      RECT 0.587 1.119 0.629 1.161 ;
      RECT 0.891 1.09 0.933 1.132 ;
      RECT 0.891 0.998 0.933 1.04 ;
      RECT 0.891 0.904 0.933 0.946 ;
      RECT 0.587 0.288 0.629 0.33 ;
      RECT 0.283 0.288 0.325 0.33 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.635 1.773 ;
  END
END NOR2X1_RVT

MACRO XNOR3X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.648 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.967 1.497 1.009 1.539 ;
      LAYER M1 ;
        RECT 0.962 1.465 1.119 1.575 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.057 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.575 0.738 1.617 0.78 ;
        RECT 0.663 0.757 0.705 0.799 ;
      LAYER M1 ;
        RECT 0.66 0.826 1.621 0.876 ;
        RECT 0.66 0.705 0.815 0.826 ;
        RECT 1.571 0.703 1.621 0.826 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0555 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 2.487 0.121 2.529 0.163 ;
        RECT 2.943 0.591 2.985 0.633 ;
      LAYER M1 ;
        RECT 2.706 0.619 2.99 0.669 ;
        RECT 2.833 0.553 2.99 0.619 ;
        RECT 2.706 0.4 2.756 0.619 ;
        RECT 2.57 0.35 2.756 0.4 ;
        RECT 2.57 0.166 2.62 0.35 ;
        RECT 2.467 0.116 2.62 0.166 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0465 ;
  END A3
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.323 0.157 3.365 0.199 ;
        RECT 3.323 0.249 3.365 0.291 ;
        RECT 3.323 0.341 3.365 0.383 ;
        RECT 3.323 0.932 3.365 0.974 ;
        RECT 3.323 1.024 3.365 1.066 ;
        RECT 3.323 1.116 3.365 1.158 ;
        RECT 3.323 1.208 3.365 1.25 ;
        RECT 3.323 1.3 3.365 1.342 ;
        RECT 3.323 1.392 3.365 1.434 ;
        RECT 3.323 1.484 3.365 1.526 ;
      LAYER M1 ;
        RECT 3.319 0.852 3.369 1.546 ;
        RECT 3.319 0.802 3.449 0.852 ;
        RECT 3.399 0.512 3.449 0.802 ;
        RECT 3.319 0.462 3.551 0.512 ;
        RECT 3.319 0.128 3.369 0.462 ;
        RECT 3.433 0.401 3.551 0.462 ;
    END
    ANTENNADIFFAREA 0.1142 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 0.981 0.325 1.023 ;
        RECT 0.283 1.073 0.325 1.115 ;
        RECT 0.283 1.165 0.325 1.207 ;
        RECT 2.107 1.25 2.149 1.292 ;
        RECT 2.867 1.253 2.909 1.295 ;
        RECT 0.283 1.257 0.325 1.299 ;
        RECT 3.171 1.3 3.213 1.342 ;
        RECT 0.587 1.325 0.629 1.367 ;
        RECT 1.043 1.325 1.085 1.367 ;
        RECT 1.651 1.325 1.693 1.367 ;
        RECT 3.171 1.392 3.213 1.434 ;
        RECT 3.171 1.484 3.213 1.526 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
        RECT 3.095 1.651 3.137 1.693 ;
        RECT 3.247 1.651 3.289 1.693 ;
        RECT 3.399 1.651 3.441 1.693 ;
        RECT 3.551 1.651 3.593 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 3.648 1.702 ;
        RECT 0.583 1.371 0.633 1.642 ;
        RECT 1.647 1.305 1.697 1.642 ;
        RECT 0.583 1.321 1.105 1.371 ;
        RECT 0.583 1.304 0.633 1.321 ;
        RECT 0.279 0.944 0.329 1.642 ;
        RECT 2.103 1.215 2.153 1.642 ;
        RECT 3.167 1.299 3.217 1.642 ;
        RECT 2.847 1.249 3.217 1.299 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 3.399 -0.021 3.441 0.021 ;
        RECT 3.551 -0.021 3.593 0.021 ;
        RECT 3.171 0.157 3.213 0.199 ;
        RECT 1.651 0.238 1.693 0.28 ;
        RECT 3.171 0.249 3.213 0.291 ;
        RECT 2.107 0.266 2.149 0.308 ;
        RECT 0.587 0.274 0.629 0.316 ;
        RECT 1.043 0.274 1.085 0.316 ;
        RECT 0.283 0.275 0.325 0.317 ;
        RECT 2.867 0.278 2.909 0.32 ;
        RECT 0.283 0.367 0.325 0.409 ;
      LAYER M1 ;
        RECT 0.279 0.391 0.581 0.441 ;
        RECT 0.531 0.32 0.581 0.391 ;
        RECT 2.847 0.274 3.217 0.324 ;
        RECT 0.531 0.27 1.105 0.32 ;
        RECT 1.631 0.234 1.785 0.284 ;
        RECT 0.279 0.03 0.329 0.391 ;
        RECT 2.103 0.03 2.153 0.343 ;
        RECT 3.167 0.03 3.217 0.274 ;
        RECT 1.735 0.03 1.785 0.234 ;
        RECT 0 -0.03 3.648 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 2.563 1.153 2.605 1.195 ;
      RECT 2.715 0.988 2.757 1.03 ;
      RECT 2.259 0.988 2.301 1.03 ;
      RECT 0.435 1.243 0.477 1.285 ;
      RECT 2.791 1.489 2.833 1.531 ;
      RECT 3.247 0.608 3.289 0.65 ;
      RECT 1.955 0.367 1.997 0.409 ;
      RECT 2.715 0.238 2.757 0.28 ;
      RECT 1.499 0.338 1.541 0.38 ;
      RECT 1.271 0.597 1.313 0.639 ;
      RECT 1.879 0.677 1.921 0.719 ;
      RECT 1.195 0.238 1.237 0.28 ;
      RECT 0.891 0.412 0.933 0.454 ;
      RECT 0.435 0.264 0.477 0.306 ;
      RECT 1.347 0.329 1.389 0.371 ;
      RECT 0.739 0.412 0.781 0.454 ;
      RECT 2.563 1.153 2.605 1.195 ;
      RECT 2.639 0.723 2.681 0.765 ;
      RECT 3.019 0.993 3.061 1.035 ;
      RECT 1.955 1.311 1.997 1.353 ;
      RECT 1.195 1.325 1.237 1.367 ;
      RECT 1.803 1.208 1.845 1.25 ;
      RECT 1.803 0.338 1.845 0.38 ;
      RECT 2.259 0.251 2.301 0.293 ;
      RECT 1.955 1.035 1.997 1.077 ;
      RECT 2.791 0.115 2.833 0.157 ;
      RECT 0.967 0.707 1.009 0.749 ;
      RECT 2.411 1.253 2.453 1.295 ;
      RECT 2.563 0.454 2.605 0.496 ;
      RECT 1.499 1.325 1.541 1.367 ;
      RECT 1.955 0.367 1.997 0.409 ;
      RECT 2.183 0.813 2.225 0.855 ;
      RECT 2.411 0.251 2.453 0.293 ;
      RECT 0.891 1.003 0.933 1.045 ;
      RECT 1.347 1.108 1.389 1.15 ;
      RECT 0.739 1.103 0.781 1.145 ;
      RECT 3.019 0.378 3.061 0.42 ;
      RECT 1.955 1.219 1.997 1.261 ;
      RECT 1.955 0.275 1.997 0.317 ;
      RECT 1.955 1.127 1.997 1.169 ;
      RECT 0.359 0.608 0.401 0.65 ;
    LAYER M1 ;
      RECT 2.711 0.111 2.853 0.161 ;
      RECT 2.711 0.161 2.761 0.3 ;
      RECT 2.999 0.989 3.09 1.039 ;
      RECT 3.04 0.769 3.09 0.989 ;
      RECT 2.604 0.719 3.09 0.769 ;
      RECT 3.04 0.424 3.09 0.719 ;
      RECT 2.999 0.374 3.09 0.424 ;
      RECT 2.543 1.149 3.207 1.199 ;
      RECT 2.834 0.872 2.884 1.149 ;
      RECT 3.157 0.654 3.207 1.149 ;
      RECT 2.395 0.822 2.884 0.872 ;
      RECT 3.157 0.604 3.309 0.654 ;
      RECT 2.395 0.5 2.445 0.822 ;
      RECT 2.395 0.45 2.625 0.5 ;
      RECT 2.238 0.984 2.777 1.034 ;
      RECT 2.295 0.297 2.345 0.984 ;
      RECT 2.239 0.247 2.473 0.297 ;
      RECT 1.479 0.334 1.865 0.384 ;
      RECT 2.687 1.485 2.853 1.535 ;
      RECT 1.359 0.375 1.409 0.434 ;
      RECT 1.326 0.325 1.409 0.375 ;
      RECT 1.951 1.165 2.001 1.377 ;
      RECT 1.327 1.104 2.001 1.115 ;
      RECT 1.951 0.859 2.001 1.104 ;
      RECT 2.006 0.484 2.056 0.809 ;
      RECT 1.359 0.434 2.056 0.484 ;
      RECT 1.951 0.244 2.001 0.434 ;
      RECT 2.358 1.165 2.408 1.249 ;
      RECT 1.951 1.154 2.408 1.165 ;
      RECT 1.327 1.115 2.408 1.154 ;
      RECT 1.951 0.809 2.245 0.859 ;
      RECT 2.687 1.299 2.737 1.485 ;
      RECT 2.358 1.249 2.737 1.299 ;
      RECT 1.175 1.321 1.561 1.371 ;
      RECT 1.418 0.534 1.925 0.584 ;
      RECT 1.875 0.584 1.925 0.754 ;
      RECT 0.947 0.703 1.468 0.753 ;
      RECT 1.418 0.584 1.468 0.703 ;
      RECT 0.549 0.999 0.953 1.049 ;
      RECT 0.549 0.591 0.888 0.641 ;
      RECT 0.838 0.458 0.888 0.591 ;
      RECT 0.838 0.408 1.236 0.458 ;
      RECT 1.186 0.458 1.236 0.593 ;
      RECT 1.186 0.593 1.35 0.643 ;
      RECT 0.549 0.641 0.599 0.999 ;
      RECT 0.431 0.153 1.241 0.203 ;
      RECT 1.191 0.203 1.241 0.3 ;
      RECT 0.431 0.203 0.481 0.341 ;
      RECT 0.431 1.204 1.865 1.254 ;
      RECT 0.431 1.254 0.481 1.32 ;
      RECT 0.434 1.099 0.801 1.149 ;
      RECT 0.434 0.491 0.785 0.541 ;
      RECT 0.735 0.377 0.785 0.491 ;
      RECT 0.434 0.654 0.484 1.099 ;
      RECT 0.339 0.604 0.484 0.654 ;
      RECT 0.434 0.541 0.484 0.604 ;
    LAYER PO ;
      RECT 2.037 0.068 2.067 1.606 ;
      RECT 2.493 0.068 2.523 1.606 ;
      RECT 2.797 0.068 2.827 1.606 ;
      RECT 2.189 0.068 2.219 1.606 ;
      RECT 2.949 0.068 2.979 1.606 ;
      RECT 2.645 0.068 2.675 1.606 ;
      RECT 3.101 0.068 3.131 1.606 ;
      RECT 3.253 0.068 3.283 1.606 ;
      RECT 3.557 0.068 3.587 1.606 ;
      RECT 3.405 0.068 3.435 1.606 ;
      RECT 2.341 0.068 2.371 1.606 ;
      RECT 1.885 0.068 1.915 1.606 ;
      RECT 1.277 0.068 1.307 1.606 ;
      RECT 0.973 0.068 1.003 1.606 ;
      RECT 1.125 0.068 1.155 1.606 ;
      RECT 1.733 0.068 1.763 1.606 ;
      RECT 0.821 0.068 0.851 1.606 ;
      RECT 0.213 0.068 0.243 1.606 ;
      RECT 0.669 0.068 0.699 1.606 ;
      RECT 0.061 0.068 0.091 1.606 ;
      RECT 1.429 0.068 1.459 1.606 ;
      RECT 0.517 0.066 0.547 1.606 ;
      RECT 1.581 0.066 1.611 1.606 ;
      RECT 0.365 0.066 0.395 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 3.763 1.781 ;
  END
END XNOR3X1_RVT

MACRO XOR2X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.967 0.613 1.009 0.655 ;
        RECT 1.271 0.675 1.313 0.717 ;
      LAYER M1 ;
        RECT 1.001 0.671 1.348 0.721 ;
        RECT 1.001 0.663 1.051 0.671 ;
        RECT 0.857 0.553 1.051 0.663 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0336 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.575 0.709 1.617 0.751 ;
        RECT 0.663 0.735 0.705 0.777 ;
      LAYER M1 ;
        RECT 0.555 0.815 1.45 0.831 ;
        RECT 0.553 0.781 1.45 0.815 ;
        RECT 0.553 0.705 0.711 0.781 ;
        RECT 1.4 0.755 1.45 0.781 ;
        RECT 1.4 0.705 1.652 0.755 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0342 ;
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 2.259 0.183 2.301 0.225 ;
        RECT 2.259 0.275 2.301 0.317 ;
        RECT 2.259 0.367 2.301 0.409 ;
        RECT 2.259 0.459 2.301 0.501 ;
        RECT 2.259 0.961 2.301 1.003 ;
        RECT 2.259 1.073 2.301 1.115 ;
        RECT 2.259 1.165 2.301 1.207 ;
        RECT 2.259 1.257 2.301 1.299 ;
        RECT 2.259 1.349 2.301 1.391 ;
        RECT 2.259 1.441 2.301 1.483 ;
      LAYER M1 ;
        RECT 2.255 0.815 2.305 1.546 ;
        RECT 2.255 0.765 2.487 0.815 ;
        RECT 2.31 0.705 2.487 0.765 ;
        RECT 2.31 0.554 2.36 0.705 ;
        RECT 2.255 0.504 2.36 0.554 ;
        RECT 2.255 0.148 2.305 0.504 ;
    END
    ANTENNADIFFAREA 0.1193 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 2.107 0.849 2.149 0.891 ;
        RECT 2.107 0.941 2.149 0.983 ;
        RECT 0.283 0.981 0.325 1.023 ;
        RECT 2.107 1.033 2.149 1.075 ;
        RECT 0.283 1.073 0.325 1.115 ;
        RECT 2.107 1.125 2.149 1.167 ;
        RECT 0.283 1.165 0.325 1.207 ;
        RECT 2.107 1.217 2.149 1.259 ;
        RECT 0.587 1.243 0.629 1.285 ;
        RECT 1.043 1.243 1.085 1.285 ;
        RECT 1.651 1.243 1.693 1.285 ;
        RECT 2.107 1.309 2.149 1.351 ;
        RECT 2.107 1.401 2.149 1.443 ;
        RECT 2.107 1.493 2.149 1.535 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 2.584 1.702 ;
        RECT 0.279 0.944 0.329 1.642 ;
        RECT 0.583 1.208 0.633 1.642 ;
        RECT 1.039 1.208 1.089 1.642 ;
        RECT 1.647 1.208 1.697 1.642 ;
        RECT 2.103 0.814 2.153 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.107 0.17 2.149 0.212 ;
        RECT 2.107 0.262 2.149 0.304 ;
        RECT 1.651 0.274 1.693 0.316 ;
        RECT 0.283 0.275 0.325 0.317 ;
        RECT 0.587 0.304 0.629 0.346 ;
        RECT 1.043 0.304 1.085 0.346 ;
        RECT 2.107 0.354 2.149 0.396 ;
        RECT 0.283 0.367 0.325 0.409 ;
      LAYER M1 ;
        RECT 0.279 0.402 0.596 0.452 ;
        RECT 0.546 0.35 0.596 0.402 ;
        RECT 0.546 0.3 1.12 0.35 ;
        RECT 1.616 0.27 1.785 0.32 ;
        RECT 2.103 0.148 2.153 0.428 ;
        RECT 1.735 0.148 1.785 0.27 ;
        RECT 1.735 0.098 2.153 0.148 ;
        RECT 0.279 0.03 0.329 0.402 ;
        RECT 2.103 0.03 2.153 0.098 ;
        RECT 0 -0.03 2.584 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.739 1.012 0.781 1.054 ;
      RECT 1.803 1.151 1.845 1.193 ;
      RECT 0.891 1.012 0.933 1.054 ;
      RECT 2.183 0.608 2.225 0.65 ;
      RECT 0.359 0.608 0.401 0.65 ;
      RECT 0.891 0.412 0.933 0.454 ;
      RECT 1.955 1.073 1.997 1.115 ;
      RECT 1.879 0.575 1.921 0.617 ;
      RECT 1.955 1.174 1.997 1.216 ;
      RECT 1.347 0.329 1.389 0.371 ;
      RECT 1.195 0.264 1.237 0.306 ;
      RECT 1.499 1.243 1.541 1.285 ;
      RECT 1.195 1.243 1.237 1.285 ;
      RECT 0.435 1.243 0.477 1.285 ;
      RECT 0.435 1.151 0.477 1.193 ;
      RECT 0.435 0.275 0.477 0.317 ;
      RECT 1.803 1.243 1.845 1.285 ;
      RECT 1.499 0.375 1.541 0.417 ;
      RECT 1.955 0.367 1.997 0.409 ;
      RECT 1.955 0.367 1.997 0.409 ;
      RECT 1.955 0.275 1.997 0.317 ;
      RECT 1.803 0.375 1.845 0.417 ;
      RECT 1.347 1.012 1.389 1.054 ;
      RECT 0.739 0.422 0.781 0.464 ;
      RECT 1.955 1.073 1.997 1.115 ;
    LAYER M1 ;
      RECT 0.403 0.519 0.785 0.569 ;
      RECT 0.403 1.008 0.801 1.058 ;
      RECT 0.735 0.402 0.785 0.519 ;
      RECT 0.324 0.604 0.453 0.654 ;
      RECT 0.403 0.569 0.453 0.604 ;
      RECT 0.403 0.654 0.453 1.008 ;
      RECT 0.431 1.108 1.849 1.158 ;
      RECT 1.799 1.158 1.849 1.32 ;
      RECT 0.431 1.158 0.481 1.32 ;
      RECT 1.17 0.571 1.956 0.621 ;
      RECT 1.113 0.89 1.752 0.94 ;
      RECT 1.702 0.621 1.752 0.89 ;
      RECT 0.871 0.408 1.22 0.458 ;
      RECT 0.871 1.008 1.163 1.058 ;
      RECT 1.17 0.458 1.22 0.571 ;
      RECT 1.113 0.94 1.163 1.008 ;
      RECT 2.006 0.604 2.26 0.654 ;
      RECT 1.343 0.294 1.393 0.471 ;
      RECT 1.343 0.471 2.056 0.521 ;
      RECT 1.951 0.704 2.056 0.754 ;
      RECT 2.006 0.654 2.056 0.704 ;
      RECT 2.006 0.521 2.056 0.604 ;
      RECT 1.951 0.24 2.001 0.471 ;
      RECT 1.951 1.058 2.001 1.315 ;
      RECT 1.312 1.008 2.001 1.058 ;
      RECT 1.951 0.754 2.001 1.008 ;
      RECT 1.16 1.239 1.576 1.289 ;
      RECT 1.464 0.371 1.88 0.421 ;
      RECT 0.431 0.153 1.241 0.203 ;
      RECT 1.191 0.203 1.241 0.326 ;
      RECT 0.431 0.203 0.481 0.352 ;
    LAYER PO ;
      RECT 1.885 0.068 1.915 1.606 ;
      RECT 1.277 0.068 1.307 1.606 ;
      RECT 0.517 0.066 0.547 1.606 ;
      RECT 1.581 0.066 1.611 1.606 ;
      RECT 2.341 0.068 2.371 1.606 ;
      RECT 2.189 0.068 2.219 1.606 ;
      RECT 0.821 0.068 0.851 1.606 ;
      RECT 0.973 0.068 1.003 1.606 ;
      RECT 2.037 0.068 2.067 1.606 ;
      RECT 1.733 0.068 1.763 1.606 ;
      RECT 1.125 0.068 1.155 1.606 ;
      RECT 1.429 0.068 1.459 1.606 ;
      RECT 0.213 0.068 0.243 1.606 ;
      RECT 0.669 0.068 0.699 1.606 ;
      RECT 0.365 0.066 0.395 1.606 ;
      RECT 0.061 0.068 0.091 1.606 ;
      RECT 2.493 0.068 2.523 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 2.699 1.781 ;
  END
END XOR2X1_RVT

MACRO AOI21X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.89 0.553 0.932 ;
      LAYER M1 ;
        RECT 0.492 0.857 0.663 0.967 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0243 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.725 0.401 0.767 ;
      LAYER M1 ;
        RECT 0.249 0.705 0.421 0.815 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0243 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.117 0.857 0.159 ;
      LAYER M1 ;
        RECT 0.705 0.097 0.877 0.207 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0228 ;
  END A3
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.499 0.134 1.541 0.176 ;
        RECT 1.499 0.226 1.541 0.268 ;
        RECT 1.499 0.318 1.541 0.36 ;
        RECT 1.499 0.41 1.541 0.452 ;
        RECT 1.499 0.848 1.541 0.89 ;
        RECT 1.499 0.94 1.541 0.982 ;
        RECT 1.499 1.032 1.541 1.074 ;
        RECT 1.499 1.124 1.541 1.166 ;
        RECT 1.499 1.216 1.541 1.258 ;
        RECT 1.499 1.308 1.541 1.35 ;
        RECT 1.499 1.4 1.541 1.442 ;
        RECT 1.499 1.492 1.541 1.534 ;
      LAYER M1 ;
        RECT 1.495 1.271 1.545 1.554 ;
        RECT 1.465 1.161 1.575 1.271 ;
        RECT 1.495 0.853 1.545 1.161 ;
        RECT 1.495 0.803 1.585 0.853 ;
        RECT 1.535 0.48 1.585 0.803 ;
        RECT 1.495 0.43 1.585 0.48 ;
        RECT 1.495 0.114 1.545 0.43 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.043 1.041 1.085 1.083 ;
        RECT 1.347 1.124 1.389 1.166 ;
        RECT 0.283 1.133 0.325 1.175 ;
        RECT 1.043 1.133 1.085 1.175 ;
        RECT 1.347 1.216 1.389 1.258 ;
        RECT 0.283 1.225 0.325 1.267 ;
        RECT 0.587 1.225 0.629 1.267 ;
        RECT 1.043 1.225 1.085 1.267 ;
        RECT 1.347 1.308 1.389 1.35 ;
        RECT 0.283 1.317 0.325 1.359 ;
        RECT 0.587 1.317 0.629 1.359 ;
        RECT 1.043 1.317 1.085 1.359 ;
        RECT 1.347 1.4 1.389 1.442 ;
        RECT 0.283 1.409 0.325 1.451 ;
        RECT 0.587 1.409 0.629 1.451 ;
        RECT 1.043 1.409 1.085 1.451 ;
        RECT 1.347 1.492 1.389 1.534 ;
        RECT 0.283 1.501 0.325 1.543 ;
        RECT 0.587 1.501 0.629 1.543 ;
        RECT 1.043 1.501 1.085 1.543 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.824 1.702 ;
        RECT 0.279 1.113 0.329 1.642 ;
        RECT 0.583 1.205 0.633 1.642 ;
        RECT 1.039 1.021 1.089 1.642 ;
        RECT 1.342 1.104 1.392 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.347 0.134 1.389 0.176 ;
        RECT 1.347 0.226 1.389 0.268 ;
        RECT 1.347 0.318 1.389 0.36 ;
        RECT 0.283 0.408 0.325 0.45 ;
        RECT 0.739 0.408 0.781 0.45 ;
        RECT 1.043 0.408 1.085 0.45 ;
        RECT 1.347 0.41 1.389 0.452 ;
        RECT 0.283 0.5 0.325 0.542 ;
        RECT 0.739 0.5 0.781 0.542 ;
        RECT 1.043 0.5 1.085 0.542 ;
      LAYER M1 ;
        RECT 0.279 0.338 0.329 0.562 ;
        RECT 0.735 0.338 0.785 0.562 ;
        RECT 0.279 0.288 0.785 0.338 ;
        RECT 1.039 0.03 1.089 0.562 ;
        RECT 1.343 0.03 1.393 0.472 ;
        RECT 0.279 0.03 0.329 0.288 ;
        RECT 0 -0.03 1.824 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.583 0.757 1.181 0.807 ;
      RECT 0.583 0.388 0.633 0.757 ;
      RECT 0.887 0.807 0.937 1.563 ;
      RECT 0.887 0.388 0.937 0.757 ;
      RECT 1.191 0.623 1.485 0.673 ;
      RECT 1.191 1.002 1.396 1.052 ;
      RECT 1.346 0.673 1.396 1.002 ;
      RECT 1.191 0.388 1.241 0.623 ;
      RECT 1.191 1.052 1.241 1.563 ;
      RECT 1.191 1.001 1.241 1.002 ;
      RECT 0.735 1.12 0.785 1.563 ;
      RECT 0.431 1.07 0.785 1.12 ;
      RECT 0.431 1.12 0.481 1.568 ;
    LAYER PO ;
      RECT 1.581 0.063 1.611 1.604 ;
      RECT 0.213 0.064 0.243 1.613 ;
      RECT 1.429 0.064 1.459 1.604 ;
      RECT 0.973 0.064 1.003 1.613 ;
      RECT 1.277 0.059 1.307 1.613 ;
      RECT 0.517 0.064 0.547 1.613 ;
      RECT 0.061 0.064 0.091 1.613 ;
      RECT 1.733 0.063 1.763 1.604 ;
      RECT 0.365 0.059 0.395 1.613 ;
      RECT 0.821 0.059 0.851 1.613 ;
      RECT 0.669 0.064 0.699 1.613 ;
      RECT 1.125 0.059 1.155 1.613 ;
    LAYER CO ;
      RECT 0.891 0.5 0.933 0.542 ;
      RECT 1.195 1.133 1.237 1.175 ;
      RECT 1.195 1.225 1.237 1.267 ;
      RECT 1.195 1.317 1.237 1.359 ;
      RECT 1.195 1.041 1.237 1.083 ;
      RECT 1.195 1.501 1.237 1.543 ;
      RECT 1.195 1.409 1.237 1.451 ;
      RECT 0.739 1.225 0.781 1.267 ;
      RECT 0.891 1.225 0.933 1.267 ;
      RECT 1.195 0.408 1.237 0.45 ;
      RECT 0.435 1.501 0.477 1.543 ;
      RECT 0.891 0.408 0.933 0.45 ;
      RECT 1.195 0.5 1.237 0.542 ;
      RECT 0.739 1.317 0.781 1.359 ;
      RECT 1.119 0.761 1.161 0.803 ;
      RECT 0.891 1.317 0.933 1.359 ;
      RECT 0.435 1.317 0.477 1.359 ;
      RECT 0.739 1.409 0.781 1.451 ;
      RECT 0.435 1.225 0.477 1.267 ;
      RECT 0.891 1.409 0.933 1.451 ;
      RECT 0.587 0.408 0.629 0.45 ;
      RECT 0.891 1.501 0.933 1.543 ;
      RECT 0.435 1.409 0.477 1.451 ;
      RECT 0.587 0.5 0.629 0.542 ;
      RECT 1.423 0.627 1.465 0.669 ;
      RECT 0.435 1.133 0.477 1.175 ;
      RECT 0.739 1.501 0.781 1.543 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.939 1.787 ;
  END
END AOI21X1_RVT

MACRO XOR3X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 4.256 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 2.335 0.596 2.377 0.638 ;
        RECT 1.119 0.615 1.161 0.657 ;
        RECT 2.487 0.677 2.529 0.719 ;
      LAYER M1 ;
        RECT 1.114 0.664 1.772 0.714 ;
        RECT 2.483 0.642 2.533 0.754 ;
        RECT 1.114 0.553 1.271 0.664 ;
        RECT 1.722 0.642 1.772 0.664 ;
        RECT 1.722 0.592 2.533 0.642 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0783 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.879 0.738 1.921 0.78 ;
        RECT 2.031 0.738 2.073 0.78 ;
        RECT 0.815 0.757 0.857 0.799 ;
      LAYER M1 ;
        RECT 0.812 0.803 2.077 0.853 ;
        RECT 0.812 0.705 0.967 0.803 ;
        RECT 1.875 0.703 1.925 0.803 ;
        RECT 2.027 0.703 2.077 0.803 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0753 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.095 0.65 3.137 0.692 ;
        RECT 3.551 0.877 3.593 0.919 ;
      LAYER M1 ;
        RECT 3.546 0.854 3.705 0.97 ;
        RECT 3.547 0.669 3.597 0.854 ;
        RECT 3.091 0.669 3.141 0.731 ;
        RECT 3.091 0.619 3.597 0.669 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0498 ;
  END A3
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.931 0.157 3.973 0.199 ;
        RECT 3.931 0.249 3.973 0.291 ;
        RECT 3.931 0.341 3.973 0.383 ;
        RECT 3.931 0.433 3.973 0.475 ;
        RECT 3.931 1.392 3.973 1.434 ;
        RECT 3.931 1.484 3.973 1.526 ;
      LAYER M1 ;
        RECT 3.927 1.299 3.977 1.546 ;
        RECT 3.927 1.249 4.057 1.299 ;
        RECT 4.007 1.119 4.057 1.249 ;
        RECT 4.007 1.009 4.159 1.119 ;
        RECT 4.007 0.542 4.057 1.009 ;
        RECT 3.927 0.492 4.057 0.542 ;
        RECT 3.927 0.127 3.977 0.492 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.435 1.243 0.477 1.285 ;
        RECT 2.715 1.25 2.757 1.292 ;
        RECT 0.739 1.253 0.781 1.295 ;
        RECT 1.195 1.253 1.237 1.295 ;
        RECT 1.955 1.253 1.997 1.295 ;
        RECT 0.435 1.335 0.477 1.377 ;
        RECT 3.475 1.361 3.517 1.403 ;
        RECT 3.779 1.401 3.821 1.443 ;
        RECT 3.779 1.493 3.821 1.535 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
        RECT 3.095 1.651 3.137 1.693 ;
        RECT 3.247 1.651 3.289 1.693 ;
        RECT 3.399 1.651 3.441 1.693 ;
        RECT 3.551 1.651 3.593 1.693 ;
        RECT 3.703 1.651 3.745 1.693 ;
        RECT 3.855 1.651 3.897 1.693 ;
        RECT 4.007 1.651 4.049 1.693 ;
        RECT 4.159 1.651 4.201 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 4.256 1.702 ;
        RECT 0.431 1.223 0.481 1.642 ;
        RECT 0.735 1.218 0.785 1.642 ;
        RECT 1.191 1.218 1.241 1.642 ;
        RECT 1.951 1.218 2.001 1.642 ;
        RECT 2.711 1.215 2.761 1.642 ;
        RECT 3.775 1.407 3.825 1.642 ;
        RECT 3.455 1.357 3.825 1.407 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 3.399 -0.021 3.441 0.021 ;
        RECT 3.551 -0.021 3.593 0.021 ;
        RECT 3.703 -0.021 3.745 0.021 ;
        RECT 3.855 -0.021 3.897 0.021 ;
        RECT 4.007 -0.021 4.049 0.021 ;
        RECT 4.159 -0.021 4.201 0.021 ;
        RECT 3.779 0.157 3.821 0.199 ;
        RECT 3.475 0.215 3.517 0.257 ;
        RECT 2.715 0.264 2.757 0.306 ;
        RECT 1.955 0.267 1.997 0.309 ;
        RECT 0.739 0.274 0.781 0.316 ;
        RECT 1.195 0.274 1.237 0.316 ;
        RECT 0.435 0.33 0.477 0.372 ;
      LAYER M1 ;
        RECT 0.162 0.391 0.733 0.441 ;
        RECT 0.683 0.32 0.733 0.391 ;
        RECT 0.431 0.3 0.481 0.391 ;
        RECT 0.683 0.27 1.272 0.32 ;
        RECT 1.92 0.263 2.241 0.313 ;
        RECT 3.45 0.211 3.843 0.261 ;
        RECT 0.162 0.03 0.212 0.391 ;
        RECT 2.711 0.03 2.761 0.326 ;
        RECT 2.191 0.03 2.241 0.263 ;
        RECT 3.775 0.03 3.825 0.211 ;
        RECT 0 -0.03 4.256 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 3.627 0.422 3.669 0.464 ;
      RECT 2.563 0.959 2.605 1.001 ;
      RECT 2.563 0.275 2.605 0.317 ;
      RECT 2.563 0.867 2.605 0.909 ;
      RECT 0.511 0.608 0.553 0.65 ;
      RECT 1.651 0.238 1.693 0.28 ;
      RECT 1.423 0.568 1.465 0.61 ;
      RECT 2.259 1.012 2.301 1.054 ;
      RECT 2.259 0.468 2.301 0.51 ;
      RECT 2.107 0.908 2.149 0.95 ;
      RECT 2.107 0.368 2.149 0.41 ;
      RECT 0.359 0.608 0.401 0.65 ;
      RECT 0.283 0.264 0.325 0.306 ;
      RECT 2.563 1.235 2.605 1.277 ;
      RECT 2.563 1.143 2.605 1.185 ;
      RECT 3.171 1.153 3.213 1.195 ;
      RECT 3.019 0.984 3.061 1.026 ;
      RECT 2.867 0.984 2.909 1.026 ;
      RECT 0.587 1.243 0.629 1.285 ;
      RECT 3.399 1.538 3.441 1.58 ;
      RECT 3.855 0.608 3.897 0.65 ;
      RECT 2.563 0.367 2.605 0.409 ;
      RECT 3.019 0.264 3.061 0.306 ;
      RECT 1.803 0.368 1.845 0.41 ;
      RECT 1.575 0.568 1.617 0.61 ;
      RECT 1.347 0.238 1.389 0.28 ;
      RECT 1.043 0.412 1.085 0.454 ;
      RECT 1.651 0.908 1.693 0.95 ;
      RECT 0.587 0.264 0.629 0.306 ;
      RECT 1.499 0.329 1.541 0.371 ;
      RECT 0.891 0.412 0.933 0.454 ;
      RECT 3.171 1.153 3.213 1.195 ;
      RECT 3.247 0.723 3.289 0.765 ;
      RECT 3.627 1.033 3.669 1.075 ;
      RECT 0.283 1.243 0.325 1.285 ;
      RECT 1.347 0.908 1.389 0.95 ;
      RECT 2.411 1.243 2.453 1.285 ;
      RECT 2.411 0.368 2.453 0.41 ;
      RECT 2.867 0.422 2.909 0.464 ;
      RECT 2.563 1.051 2.605 1.093 ;
      RECT 3.399 0.115 3.441 0.157 ;
      RECT 3.323 1.253 3.365 1.295 ;
      RECT 3.171 0.322 3.213 0.364 ;
      RECT 1.803 0.908 1.845 0.95 ;
      RECT 2.563 0.367 2.605 0.409 ;
      RECT 2.791 0.608 2.833 0.65 ;
      RECT 3.323 0.422 3.365 0.464 ;
      RECT 1.043 0.985 1.085 1.027 ;
      RECT 1.499 1.012 1.541 1.054 ;
      RECT 0.891 1.022 0.933 1.064 ;
    LAYER M1 ;
      RECT 3.321 1.534 3.461 1.584 ;
      RECT 1.479 0.325 1.58 0.375 ;
      RECT 1.53 0.375 1.58 0.464 ;
      RECT 1.53 0.464 2.664 0.514 ;
      RECT 2.559 1.165 2.609 1.305 ;
      RECT 2.559 0.809 2.664 0.859 ;
      RECT 2.559 1.058 2.609 1.115 ;
      RECT 1.464 1.008 2.609 1.058 ;
      RECT 2.614 0.654 2.664 0.809 ;
      RECT 2.559 0.241 2.609 0.464 ;
      RECT 2.614 0.514 2.664 0.604 ;
      RECT 2.559 0.859 2.609 1.008 ;
      RECT 3.007 1.249 3.385 1.299 ;
      RECT 3.321 1.299 3.371 1.534 ;
      RECT 3.007 1.165 3.057 1.249 ;
      RECT 2.559 1.115 3.057 1.165 ;
      RECT 2.787 0.654 2.837 0.685 ;
      RECT 2.787 0.573 2.837 0.604 ;
      RECT 2.614 0.604 2.837 0.654 ;
      RECT 0.397 1.018 0.953 1.068 ;
      RECT 0.397 0.491 0.937 0.541 ;
      RECT 0.887 0.377 0.937 0.491 ;
      RECT 0.339 0.604 0.573 0.654 ;
      RECT 0.397 0.541 0.447 0.604 ;
      RECT 0.397 0.654 0.447 1.018 ;
      RECT 0.999 0.408 1.408 0.458 ;
      RECT 1.358 0.458 1.408 0.564 ;
      RECT 1.358 0.564 1.654 0.614 ;
      RECT 0.632 0.918 1.089 0.968 ;
      RECT 1.039 0.968 1.089 1.068 ;
      RECT 0.632 0.591 1.049 0.641 ;
      RECT 0.999 0.458 1.049 0.591 ;
      RECT 0.632 0.641 0.682 0.918 ;
      RECT 0.279 0.153 1.697 0.203 ;
      RECT 1.343 0.203 1.393 0.3 ;
      RECT 1.647 0.203 1.697 0.3 ;
      RECT 0.279 0.203 0.329 0.341 ;
      RECT 0.583 0.203 0.633 0.341 ;
      RECT 3.592 0.418 3.745 0.468 ;
      RECT 3.298 1.029 3.822 1.079 ;
      RECT 3.695 0.468 3.745 0.71 ;
      RECT 3.695 0.71 3.822 0.76 ;
      RECT 3.772 0.76 3.822 1.029 ;
      RECT 3.298 0.769 3.348 1.029 ;
      RECT 3.212 0.719 3.348 0.769 ;
      RECT 1.783 0.364 2.488 0.414 ;
      RECT 3.821 0.604 3.932 0.654 ;
      RECT 3.15 1.149 3.931 1.199 ;
      RECT 3.881 0.654 3.931 1.149 ;
      RECT 2.987 0.569 3.037 0.822 ;
      RECT 2.987 0.822 3.23 0.872 ;
      RECT 2.987 0.519 3.485 0.569 ;
      RECT 3.435 0.368 3.485 0.519 ;
      RECT 3.131 0.318 3.485 0.368 ;
      RECT 3.18 0.872 3.23 1.149 ;
      RECT 0.279 1.118 2.457 1.168 ;
      RECT 2.407 1.168 2.457 1.32 ;
      RECT 0.279 1.168 0.329 1.32 ;
      RECT 0.583 1.168 0.633 1.32 ;
      RECT 3.015 0.111 3.461 0.161 ;
      RECT 3.015 0.161 3.065 0.326 ;
      RECT 2.827 0.98 3.096 1.03 ;
      RECT 2.847 0.418 3.385 0.468 ;
      RECT 2.887 0.468 2.937 0.98 ;
      RECT 1.327 0.904 2.169 0.954 ;
    LAYER PO ;
      RECT 1.429 0.068 1.459 1.606 ;
      RECT 1.581 0.068 1.611 1.606 ;
      RECT 2.493 0.068 2.523 1.606 ;
      RECT 2.341 0.068 2.371 1.606 ;
      RECT 1.885 0.066 1.915 1.606 ;
      RECT 2.037 0.066 2.067 1.606 ;
      RECT 0.365 0.066 0.395 1.606 ;
      RECT 2.645 0.068 2.675 1.606 ;
      RECT 3.101 0.068 3.131 1.606 ;
      RECT 3.405 0.068 3.435 1.606 ;
      RECT 2.797 0.068 2.827 1.606 ;
      RECT 3.557 0.068 3.587 1.606 ;
      RECT 3.253 0.068 3.283 1.606 ;
      RECT 3.709 0.068 3.739 1.606 ;
      RECT 3.861 0.068 3.891 1.606 ;
      RECT 4.165 0.068 4.195 1.606 ;
      RECT 4.013 0.068 4.043 1.606 ;
      RECT 2.949 0.068 2.979 1.606 ;
      RECT 0.517 0.066 0.547 1.606 ;
      RECT 1.125 0.068 1.155 1.606 ;
      RECT 1.277 0.068 1.307 1.606 ;
      RECT 2.189 0.068 2.219 1.606 ;
      RECT 0.973 0.068 1.003 1.606 ;
      RECT 0.213 0.068 0.243 1.606 ;
      RECT 0.821 0.068 0.851 1.606 ;
      RECT 0.061 0.068 0.091 1.606 ;
      RECT 1.733 0.068 1.763 1.606 ;
      RECT 0.669 0.066 0.699 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 4.371 1.773 ;
  END
END XOR3X1_RVT

MACRO AO221X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.893 0.401 0.935 ;
      LAYER M1 ;
        RECT 0.249 0.857 0.404 0.967 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0249 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.607 0.553 0.649 ;
      LAYER M1 ;
        RECT 0.401 0.553 0.573 0.663 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0249 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.132 0.857 0.174 ;
      LAYER M1 ;
        RECT 0.705 0.097 0.863 0.207 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0249 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.896 0.705 0.938 ;
      LAYER M1 ;
        RECT 0.553 1.009 0.663 1.119 ;
        RECT 0.613 0.942 0.663 1.009 ;
        RECT 0.613 0.893 0.725 0.942 ;
        RECT 0.623 0.892 0.725 0.893 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0249 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.119 0.777 1.161 0.819 ;
      LAYER M1 ;
        RECT 1.009 0.773 1.181 0.823 ;
        RECT 1.009 0.705 1.119 0.773 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.021 ;
  END A5
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.499 0.166 1.541 0.208 ;
        RECT 1.499 0.258 1.541 0.3 ;
        RECT 1.499 0.35 1.541 0.392 ;
        RECT 1.499 0.442 1.541 0.484 ;
        RECT 1.499 0.86 1.541 0.902 ;
        RECT 1.499 0.952 1.541 0.994 ;
        RECT 1.499 1.044 1.541 1.086 ;
        RECT 1.499 1.136 1.541 1.178 ;
        RECT 1.499 1.228 1.541 1.27 ;
        RECT 1.499 1.32 1.541 1.362 ;
        RECT 1.499 1.412 1.541 1.454 ;
        RECT 1.499 1.504 1.541 1.546 ;
      LAYER M1 ;
        RECT 1.495 1.271 1.545 1.566 ;
        RECT 1.465 1.161 1.575 1.271 ;
        RECT 1.495 0.865 1.545 1.161 ;
        RECT 1.495 0.864 1.585 0.865 ;
        RECT 1.495 0.815 1.595 0.864 ;
        RECT 1.545 0.504 1.595 0.815 ;
        RECT 1.495 0.453 1.595 0.504 ;
        RECT 1.495 0.146 1.545 0.453 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.347 0.768 1.389 0.81 ;
        RECT 1.347 0.86 1.389 0.902 ;
        RECT 1.347 0.952 1.389 0.994 ;
        RECT 1.347 1.044 1.389 1.086 ;
        RECT 1.347 1.136 1.389 1.178 ;
        RECT 1.347 1.228 1.389 1.27 ;
        RECT 1.347 1.32 1.389 1.362 ;
        RECT 0.435 1.407 0.477 1.449 ;
        RECT 1.347 1.412 1.389 1.454 ;
        RECT 0.435 1.499 0.477 1.541 ;
        RECT 1.347 1.504 1.389 1.546 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.824 1.702 ;
        RECT 0.431 1.387 0.481 1.642 ;
        RECT 1.342 0.748 1.392 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.347 0.146 1.389 0.188 ;
        RECT 1.347 0.238 1.389 0.28 ;
        RECT 1.043 0.304 1.085 0.346 ;
        RECT 0.587 0.317 0.629 0.359 ;
        RECT 1.347 0.33 1.389 0.372 ;
        RECT 0.587 0.409 0.629 0.451 ;
        RECT 1.347 0.422 1.389 0.464 ;
      LAYER M1 ;
        RECT 1.343 0.03 1.393 0.484 ;
        RECT 0.583 0.03 0.633 0.471 ;
        RECT 1.04 0.03 1.09 0.366 ;
        RECT 0 -0.03 1.824 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.191 0.635 1.485 0.685 ;
      RECT 0.279 0.296 0.329 0.728 ;
      RECT 0.279 0.728 0.937 0.778 ;
      RECT 0.887 0.778 0.937 0.908 ;
      RECT 0.887 0.56 0.937 0.728 ;
      RECT 0.887 0.321 0.937 0.51 ;
      RECT 1.191 0.958 1.241 1.571 ;
      RECT 0.887 0.908 1.241 0.958 ;
      RECT 1.191 0.56 1.241 0.635 ;
      RECT 1.191 0.266 1.241 0.51 ;
      RECT 0.887 0.51 1.241 0.56 ;
      RECT 0.887 1.337 0.937 1.57 ;
      RECT 0.583 1.337 0.633 1.57 ;
      RECT 0.279 1.287 0.937 1.337 ;
      RECT 0.279 1.337 0.329 1.57 ;
      RECT 1.039 1.071 1.089 1.571 ;
      RECT 0.735 1.021 1.089 1.071 ;
      RECT 0.735 1.071 0.785 1.237 ;
    LAYER PO ;
      RECT 1.277 0.075 1.307 1.616 ;
      RECT 1.581 0.075 1.611 1.616 ;
      RECT 1.125 0.076 1.155 1.621 ;
      RECT 0.213 0.072 0.243 1.621 ;
      RECT 0.821 0.072 0.851 1.621 ;
      RECT 1.429 0.076 1.459 1.616 ;
      RECT 0.973 0.076 1.003 1.621 ;
      RECT 0.061 0.072 0.091 1.621 ;
      RECT 1.733 0.075 1.763 1.616 ;
      RECT 0.365 0.067 0.395 1.621 ;
      RECT 0.517 0.072 0.547 1.621 ;
      RECT 0.669 0.072 0.699 1.621 ;
    LAYER CO ;
      RECT 0.891 1.508 0.933 1.55 ;
      RECT 0.891 0.341 0.933 0.383 ;
      RECT 0.891 1.416 0.933 1.458 ;
      RECT 1.423 0.639 1.465 0.681 ;
      RECT 0.891 0.433 0.933 0.475 ;
      RECT 0.283 0.408 0.325 0.45 ;
      RECT 0.587 1.324 0.629 1.366 ;
      RECT 0.587 1.416 0.629 1.458 ;
      RECT 0.739 1.083 0.781 1.125 ;
      RECT 0.739 1.175 0.781 1.217 ;
      RECT 0.283 1.508 0.325 1.55 ;
      RECT 0.283 1.416 0.325 1.458 ;
      RECT 0.891 1.324 0.933 1.366 ;
      RECT 0.283 1.324 0.325 1.366 ;
      RECT 0.587 1.508 0.629 1.55 ;
      RECT 1.043 1.233 1.085 1.275 ;
      RECT 1.043 1.417 1.085 1.459 ;
      RECT 1.043 1.325 1.085 1.367 ;
      RECT 1.195 0.304 1.237 0.346 ;
      RECT 1.043 1.509 1.085 1.551 ;
      RECT 1.195 1.509 1.237 1.551 ;
      RECT 1.195 1.141 1.237 1.183 ;
      RECT 1.195 1.233 1.237 1.275 ;
      RECT 1.195 1.417 1.237 1.459 ;
      RECT 1.195 1.325 1.237 1.367 ;
      RECT 1.043 1.141 1.085 1.183 ;
      RECT 1.195 1.049 1.237 1.091 ;
      RECT 1.043 1.049 1.085 1.091 ;
      RECT 0.283 0.316 0.325 0.358 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.939 1.773 ;
  END
END AO221X1_RVT

MACRO INVX32_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 5.472 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.664 0.401 0.706 ;
        RECT 0.511 0.664 0.553 0.706 ;
        RECT 0.663 0.664 0.705 0.706 ;
        RECT 0.815 0.664 0.857 0.706 ;
        RECT 0.967 0.664 1.009 0.706 ;
        RECT 1.119 0.664 1.161 0.706 ;
        RECT 1.271 0.664 1.313 0.706 ;
        RECT 1.423 0.664 1.465 0.706 ;
        RECT 1.575 0.664 1.617 0.706 ;
        RECT 1.727 0.664 1.769 0.706 ;
        RECT 1.879 0.664 1.921 0.706 ;
        RECT 2.031 0.664 2.073 0.706 ;
        RECT 2.183 0.664 2.225 0.706 ;
        RECT 2.335 0.664 2.377 0.706 ;
        RECT 2.487 0.664 2.529 0.706 ;
        RECT 2.639 0.664 2.681 0.706 ;
        RECT 2.791 0.664 2.833 0.706 ;
        RECT 2.943 0.664 2.985 0.706 ;
        RECT 3.095 0.664 3.137 0.706 ;
        RECT 3.247 0.664 3.289 0.706 ;
        RECT 3.399 0.664 3.441 0.706 ;
        RECT 3.551 0.664 3.593 0.706 ;
        RECT 3.703 0.664 3.745 0.706 ;
        RECT 3.855 0.664 3.897 0.706 ;
        RECT 4.007 0.664 4.049 0.706 ;
        RECT 4.159 0.664 4.201 0.706 ;
        RECT 4.311 0.664 4.353 0.706 ;
        RECT 4.463 0.664 4.505 0.706 ;
        RECT 4.615 0.664 4.657 0.706 ;
        RECT 4.767 0.664 4.809 0.706 ;
        RECT 4.919 0.664 4.961 0.706 ;
        RECT 5.071 0.664 5.113 0.706 ;
      LAYER M1 ;
        RECT 0.249 0.71 0.362 0.815 ;
        RECT 0.249 0.66 5.148 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1712 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.283 0.151 0.325 0.193 ;
        RECT 0.587 0.151 0.629 0.193 ;
        RECT 0.891 0.151 0.933 0.193 ;
        RECT 1.195 0.151 1.237 0.193 ;
        RECT 1.803 0.151 1.845 0.193 ;
        RECT 2.107 0.151 2.149 0.193 ;
        RECT 2.411 0.151 2.453 0.193 ;
        RECT 2.715 0.151 2.757 0.193 ;
        RECT 3.019 0.151 3.061 0.193 ;
        RECT 3.323 0.151 3.365 0.193 ;
        RECT 3.627 0.151 3.669 0.193 ;
        RECT 3.931 0.151 3.973 0.193 ;
        RECT 4.235 0.151 4.277 0.193 ;
        RECT 4.539 0.151 4.581 0.193 ;
        RECT 4.843 0.151 4.885 0.193 ;
        RECT 5.147 0.151 5.189 0.193 ;
        RECT 1.499 0.152 1.541 0.194 ;
        RECT 0.283 0.243 0.325 0.285 ;
        RECT 0.587 0.243 0.629 0.285 ;
        RECT 0.891 0.243 0.933 0.285 ;
        RECT 1.195 0.243 1.237 0.285 ;
        RECT 1.803 0.243 1.845 0.285 ;
        RECT 2.107 0.243 2.149 0.285 ;
        RECT 2.411 0.243 2.453 0.285 ;
        RECT 2.715 0.243 2.757 0.285 ;
        RECT 3.019 0.243 3.061 0.285 ;
        RECT 3.323 0.243 3.365 0.285 ;
        RECT 3.627 0.243 3.669 0.285 ;
        RECT 3.931 0.243 3.973 0.285 ;
        RECT 4.235 0.243 4.277 0.285 ;
        RECT 4.539 0.243 4.581 0.285 ;
        RECT 4.843 0.243 4.885 0.285 ;
        RECT 5.147 0.243 5.189 0.285 ;
        RECT 1.499 0.244 1.541 0.286 ;
        RECT 0.283 0.335 0.325 0.377 ;
        RECT 0.587 0.335 0.629 0.377 ;
        RECT 0.891 0.335 0.933 0.377 ;
        RECT 1.195 0.335 1.237 0.377 ;
        RECT 1.803 0.335 1.845 0.377 ;
        RECT 2.107 0.335 2.149 0.377 ;
        RECT 2.411 0.335 2.453 0.377 ;
        RECT 2.715 0.335 2.757 0.377 ;
        RECT 3.019 0.335 3.061 0.377 ;
        RECT 3.323 0.335 3.365 0.377 ;
        RECT 3.627 0.335 3.669 0.377 ;
        RECT 3.931 0.335 3.973 0.377 ;
        RECT 4.235 0.335 4.277 0.377 ;
        RECT 4.539 0.335 4.581 0.377 ;
        RECT 4.843 0.335 4.885 0.377 ;
        RECT 5.147 0.335 5.189 0.377 ;
        RECT 1.499 0.336 1.541 0.378 ;
        RECT 0.283 0.427 0.325 0.469 ;
        RECT 0.587 0.427 0.629 0.469 ;
        RECT 0.891 0.427 0.933 0.469 ;
        RECT 1.195 0.427 1.237 0.469 ;
        RECT 1.803 0.427 1.845 0.469 ;
        RECT 2.107 0.427 2.149 0.469 ;
        RECT 2.411 0.427 2.453 0.469 ;
        RECT 2.715 0.427 2.757 0.469 ;
        RECT 3.019 0.427 3.061 0.469 ;
        RECT 3.323 0.427 3.365 0.469 ;
        RECT 3.627 0.427 3.669 0.469 ;
        RECT 3.931 0.427 3.973 0.469 ;
        RECT 4.235 0.427 4.277 0.469 ;
        RECT 4.539 0.427 4.581 0.469 ;
        RECT 4.843 0.427 4.885 0.469 ;
        RECT 5.147 0.427 5.189 0.469 ;
        RECT 1.499 0.428 1.541 0.47 ;
        RECT 0.283 1.027 0.325 1.069 ;
        RECT 0.587 1.027 0.629 1.069 ;
        RECT 0.891 1.027 0.933 1.069 ;
        RECT 1.195 1.027 1.237 1.069 ;
        RECT 1.803 1.027 1.845 1.069 ;
        RECT 2.107 1.027 2.149 1.069 ;
        RECT 2.411 1.027 2.453 1.069 ;
        RECT 2.715 1.027 2.757 1.069 ;
        RECT 3.019 1.027 3.061 1.069 ;
        RECT 3.323 1.027 3.365 1.069 ;
        RECT 3.627 1.027 3.669 1.069 ;
        RECT 3.931 1.027 3.973 1.069 ;
        RECT 4.235 1.027 4.277 1.069 ;
        RECT 4.539 1.027 4.581 1.069 ;
        RECT 4.843 1.027 4.885 1.069 ;
        RECT 5.147 1.027 5.189 1.069 ;
        RECT 1.499 1.028 1.541 1.07 ;
        RECT 0.283 1.119 0.325 1.161 ;
        RECT 0.587 1.119 0.629 1.161 ;
        RECT 0.891 1.119 0.933 1.161 ;
        RECT 1.195 1.119 1.237 1.161 ;
        RECT 1.803 1.119 1.845 1.161 ;
        RECT 2.107 1.119 2.149 1.161 ;
        RECT 2.411 1.119 2.453 1.161 ;
        RECT 2.715 1.119 2.757 1.161 ;
        RECT 3.019 1.119 3.061 1.161 ;
        RECT 3.323 1.119 3.365 1.161 ;
        RECT 3.627 1.119 3.669 1.161 ;
        RECT 3.931 1.119 3.973 1.161 ;
        RECT 4.235 1.119 4.277 1.161 ;
        RECT 4.539 1.119 4.581 1.161 ;
        RECT 4.843 1.119 4.885 1.161 ;
        RECT 5.147 1.119 5.189 1.161 ;
        RECT 1.499 1.12 1.541 1.162 ;
        RECT 0.283 1.211 0.325 1.253 ;
        RECT 0.587 1.211 0.629 1.253 ;
        RECT 0.891 1.211 0.933 1.253 ;
        RECT 1.195 1.211 1.237 1.253 ;
        RECT 1.803 1.211 1.845 1.253 ;
        RECT 2.107 1.211 2.149 1.253 ;
        RECT 2.411 1.211 2.453 1.253 ;
        RECT 2.715 1.211 2.757 1.253 ;
        RECT 3.019 1.211 3.061 1.253 ;
        RECT 3.323 1.211 3.365 1.253 ;
        RECT 3.627 1.211 3.669 1.253 ;
        RECT 3.931 1.211 3.973 1.253 ;
        RECT 4.235 1.211 4.277 1.253 ;
        RECT 4.539 1.211 4.581 1.253 ;
        RECT 4.843 1.211 4.885 1.253 ;
        RECT 5.147 1.211 5.189 1.253 ;
        RECT 1.499 1.212 1.541 1.254 ;
        RECT 0.283 1.303 0.325 1.345 ;
        RECT 0.587 1.303 0.629 1.345 ;
        RECT 0.891 1.303 0.933 1.345 ;
        RECT 1.195 1.303 1.237 1.345 ;
        RECT 1.803 1.303 1.845 1.345 ;
        RECT 2.107 1.303 2.149 1.345 ;
        RECT 2.411 1.303 2.453 1.345 ;
        RECT 2.715 1.303 2.757 1.345 ;
        RECT 3.019 1.303 3.061 1.345 ;
        RECT 3.323 1.303 3.365 1.345 ;
        RECT 3.627 1.303 3.669 1.345 ;
        RECT 3.931 1.303 3.973 1.345 ;
        RECT 4.235 1.303 4.277 1.345 ;
        RECT 4.539 1.303 4.581 1.345 ;
        RECT 4.843 1.303 4.885 1.345 ;
        RECT 5.147 1.303 5.189 1.345 ;
        RECT 1.499 1.304 1.541 1.346 ;
        RECT 0.283 1.395 0.325 1.437 ;
        RECT 0.587 1.395 0.629 1.437 ;
        RECT 0.891 1.395 0.933 1.437 ;
        RECT 1.195 1.395 1.237 1.437 ;
        RECT 1.803 1.395 1.845 1.437 ;
        RECT 2.107 1.395 2.149 1.437 ;
        RECT 2.411 1.395 2.453 1.437 ;
        RECT 2.715 1.395 2.757 1.437 ;
        RECT 3.019 1.395 3.061 1.437 ;
        RECT 3.323 1.395 3.365 1.437 ;
        RECT 3.627 1.395 3.669 1.437 ;
        RECT 3.931 1.395 3.973 1.437 ;
        RECT 4.235 1.395 4.277 1.437 ;
        RECT 4.539 1.395 4.581 1.437 ;
        RECT 4.843 1.395 4.885 1.437 ;
        RECT 5.147 1.395 5.189 1.437 ;
        RECT 1.499 1.396 1.541 1.438 ;
        RECT 0.283 1.487 0.325 1.529 ;
        RECT 0.587 1.487 0.629 1.529 ;
        RECT 0.891 1.487 0.933 1.529 ;
        RECT 1.195 1.487 1.237 1.529 ;
        RECT 1.803 1.487 1.845 1.529 ;
        RECT 2.107 1.487 2.149 1.529 ;
        RECT 2.411 1.487 2.453 1.529 ;
        RECT 2.715 1.487 2.757 1.529 ;
        RECT 3.019 1.487 3.061 1.529 ;
        RECT 3.323 1.487 3.365 1.529 ;
        RECT 3.627 1.487 3.669 1.529 ;
        RECT 3.931 1.487 3.973 1.529 ;
        RECT 4.235 1.487 4.277 1.529 ;
        RECT 4.539 1.487 4.581 1.529 ;
        RECT 4.843 1.487 4.885 1.529 ;
        RECT 5.147 1.487 5.189 1.529 ;
        RECT 1.499 1.488 1.541 1.53 ;
      LAYER M1 ;
        RECT 3.015 0.942 3.065 1.564 ;
        RECT 3.319 0.942 3.369 1.564 ;
        RECT 3.623 0.942 3.673 1.564 ;
        RECT 3.927 0.942 3.977 1.564 ;
        RECT 4.231 0.942 4.281 1.564 ;
        RECT 4.535 0.942 4.585 1.564 ;
        RECT 4.839 0.942 4.889 1.564 ;
        RECT 5.143 0.942 5.193 1.564 ;
        RECT 5.202 0.663 5.252 0.892 ;
        RECT 0.279 0.892 5.252 0.942 ;
        RECT 1.495 0.942 1.545 1.565 ;
        RECT 0.279 0.942 0.329 1.564 ;
        RECT 0.583 0.942 0.633 1.564 ;
        RECT 0.887 0.942 0.937 1.564 ;
        RECT 1.191 0.942 1.241 1.564 ;
        RECT 1.799 0.942 1.849 1.564 ;
        RECT 2.103 0.942 2.153 1.564 ;
        RECT 2.407 0.942 2.457 1.564 ;
        RECT 2.711 0.942 2.761 1.564 ;
        RECT 5.202 0.587 5.375 0.663 ;
        RECT 0.279 0.537 5.375 0.587 ;
        RECT 3.015 0.116 3.065 0.537 ;
        RECT 3.319 0.116 3.369 0.537 ;
        RECT 3.623 0.116 3.673 0.537 ;
        RECT 3.927 0.116 3.977 0.537 ;
        RECT 4.231 0.116 4.281 0.537 ;
        RECT 4.535 0.116 4.585 0.537 ;
        RECT 4.839 0.116 4.889 0.537 ;
        RECT 5.143 0.116 5.193 0.537 ;
        RECT 0.279 0.116 0.329 0.537 ;
        RECT 0.583 0.116 0.633 0.537 ;
        RECT 0.887 0.116 0.937 0.537 ;
        RECT 1.191 0.116 1.241 0.537 ;
        RECT 1.495 0.117 1.545 0.537 ;
        RECT 1.799 0.116 1.849 0.537 ;
        RECT 2.103 0.116 2.153 0.537 ;
        RECT 2.407 0.116 2.457 0.537 ;
        RECT 2.711 0.116 2.761 0.537 ;
    END
    ANTENNADIFFAREA 2.4808 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.435 1.027 0.477 1.069 ;
        RECT 0.739 1.027 0.781 1.069 ;
        RECT 1.043 1.027 1.085 1.069 ;
        RECT 1.347 1.027 1.389 1.069 ;
        RECT 1.651 1.027 1.693 1.069 ;
        RECT 1.955 1.027 1.997 1.069 ;
        RECT 2.259 1.027 2.301 1.069 ;
        RECT 2.563 1.027 2.605 1.069 ;
        RECT 2.867 1.027 2.909 1.069 ;
        RECT 3.171 1.027 3.213 1.069 ;
        RECT 3.475 1.027 3.517 1.069 ;
        RECT 3.779 1.027 3.821 1.069 ;
        RECT 4.083 1.027 4.125 1.069 ;
        RECT 4.387 1.027 4.429 1.069 ;
        RECT 4.691 1.027 4.733 1.069 ;
        RECT 4.995 1.027 5.037 1.069 ;
        RECT 0.435 1.119 0.477 1.161 ;
        RECT 0.739 1.119 0.781 1.161 ;
        RECT 1.043 1.119 1.085 1.161 ;
        RECT 1.347 1.119 1.389 1.161 ;
        RECT 1.651 1.119 1.693 1.161 ;
        RECT 1.955 1.119 1.997 1.161 ;
        RECT 2.259 1.119 2.301 1.161 ;
        RECT 2.563 1.119 2.605 1.161 ;
        RECT 2.867 1.119 2.909 1.161 ;
        RECT 3.171 1.119 3.213 1.161 ;
        RECT 3.475 1.119 3.517 1.161 ;
        RECT 3.779 1.119 3.821 1.161 ;
        RECT 4.083 1.119 4.125 1.161 ;
        RECT 4.387 1.119 4.429 1.161 ;
        RECT 4.691 1.119 4.733 1.161 ;
        RECT 4.995 1.119 5.037 1.161 ;
        RECT 0.435 1.211 0.477 1.253 ;
        RECT 0.739 1.211 0.781 1.253 ;
        RECT 1.043 1.211 1.085 1.253 ;
        RECT 1.347 1.211 1.389 1.253 ;
        RECT 1.651 1.211 1.693 1.253 ;
        RECT 1.955 1.211 1.997 1.253 ;
        RECT 2.259 1.211 2.301 1.253 ;
        RECT 2.563 1.211 2.605 1.253 ;
        RECT 2.867 1.211 2.909 1.253 ;
        RECT 3.171 1.211 3.213 1.253 ;
        RECT 3.475 1.211 3.517 1.253 ;
        RECT 3.779 1.211 3.821 1.253 ;
        RECT 4.083 1.211 4.125 1.253 ;
        RECT 4.387 1.211 4.429 1.253 ;
        RECT 4.691 1.211 4.733 1.253 ;
        RECT 4.995 1.211 5.037 1.253 ;
        RECT 0.435 1.303 0.477 1.345 ;
        RECT 0.739 1.303 0.781 1.345 ;
        RECT 1.043 1.303 1.085 1.345 ;
        RECT 1.347 1.303 1.389 1.345 ;
        RECT 1.651 1.303 1.693 1.345 ;
        RECT 1.955 1.303 1.997 1.345 ;
        RECT 2.259 1.303 2.301 1.345 ;
        RECT 2.563 1.303 2.605 1.345 ;
        RECT 2.867 1.303 2.909 1.345 ;
        RECT 3.171 1.303 3.213 1.345 ;
        RECT 3.475 1.303 3.517 1.345 ;
        RECT 3.779 1.303 3.821 1.345 ;
        RECT 4.083 1.303 4.125 1.345 ;
        RECT 4.387 1.303 4.429 1.345 ;
        RECT 4.691 1.303 4.733 1.345 ;
        RECT 4.995 1.303 5.037 1.345 ;
        RECT 0.435 1.395 0.477 1.437 ;
        RECT 0.739 1.395 0.781 1.437 ;
        RECT 1.043 1.395 1.085 1.437 ;
        RECT 1.347 1.395 1.389 1.437 ;
        RECT 1.651 1.395 1.693 1.437 ;
        RECT 1.955 1.395 1.997 1.437 ;
        RECT 2.259 1.395 2.301 1.437 ;
        RECT 2.563 1.395 2.605 1.437 ;
        RECT 2.867 1.395 2.909 1.437 ;
        RECT 3.171 1.395 3.213 1.437 ;
        RECT 3.475 1.395 3.517 1.437 ;
        RECT 3.779 1.395 3.821 1.437 ;
        RECT 4.083 1.395 4.125 1.437 ;
        RECT 4.387 1.395 4.429 1.437 ;
        RECT 4.691 1.395 4.733 1.437 ;
        RECT 4.995 1.395 5.037 1.437 ;
        RECT 0.435 1.487 0.477 1.529 ;
        RECT 0.739 1.487 0.781 1.529 ;
        RECT 1.043 1.487 1.085 1.529 ;
        RECT 1.347 1.487 1.389 1.529 ;
        RECT 1.651 1.487 1.693 1.529 ;
        RECT 1.955 1.487 1.997 1.529 ;
        RECT 2.259 1.487 2.301 1.529 ;
        RECT 2.563 1.487 2.605 1.529 ;
        RECT 2.867 1.487 2.909 1.529 ;
        RECT 3.171 1.487 3.213 1.529 ;
        RECT 3.475 1.487 3.517 1.529 ;
        RECT 3.779 1.487 3.821 1.529 ;
        RECT 4.083 1.487 4.125 1.529 ;
        RECT 4.387 1.487 4.429 1.529 ;
        RECT 4.691 1.487 4.733 1.529 ;
        RECT 4.995 1.487 5.037 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
        RECT 3.095 1.651 3.137 1.693 ;
        RECT 3.247 1.651 3.289 1.693 ;
        RECT 3.399 1.651 3.441 1.693 ;
        RECT 3.551 1.651 3.593 1.693 ;
        RECT 3.703 1.651 3.745 1.693 ;
        RECT 3.855 1.651 3.897 1.693 ;
        RECT 4.007 1.651 4.049 1.693 ;
        RECT 4.159 1.651 4.201 1.693 ;
        RECT 4.311 1.651 4.353 1.693 ;
        RECT 4.463 1.651 4.505 1.693 ;
        RECT 4.615 1.651 4.657 1.693 ;
        RECT 4.767 1.651 4.809 1.693 ;
        RECT 4.919 1.651 4.961 1.693 ;
        RECT 5.071 1.651 5.113 1.693 ;
        RECT 5.223 1.651 5.265 1.693 ;
        RECT 5.375 1.651 5.417 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 5.472 1.702 ;
        RECT 2.863 0.992 2.913 1.642 ;
        RECT 3.167 0.992 3.217 1.642 ;
        RECT 3.471 0.992 3.521 1.642 ;
        RECT 3.775 0.992 3.825 1.642 ;
        RECT 4.079 0.992 4.129 1.642 ;
        RECT 4.383 0.992 4.433 1.642 ;
        RECT 4.687 0.992 4.737 1.642 ;
        RECT 4.991 0.992 5.041 1.642 ;
        RECT 0.431 0.992 0.481 1.642 ;
        RECT 0.735 0.992 0.785 1.642 ;
        RECT 1.039 0.992 1.089 1.642 ;
        RECT 1.343 0.992 1.393 1.642 ;
        RECT 1.647 0.992 1.697 1.642 ;
        RECT 1.951 0.992 2.001 1.642 ;
        RECT 2.255 0.992 2.305 1.642 ;
        RECT 2.559 0.992 2.609 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 3.399 -0.021 3.441 0.021 ;
        RECT 3.551 -0.021 3.593 0.021 ;
        RECT 3.703 -0.021 3.745 0.021 ;
        RECT 3.855 -0.021 3.897 0.021 ;
        RECT 4.007 -0.021 4.049 0.021 ;
        RECT 4.159 -0.021 4.201 0.021 ;
        RECT 4.311 -0.021 4.353 0.021 ;
        RECT 4.463 -0.021 4.505 0.021 ;
        RECT 4.615 -0.021 4.657 0.021 ;
        RECT 4.767 -0.021 4.809 0.021 ;
        RECT 4.919 -0.021 4.961 0.021 ;
        RECT 5.071 -0.021 5.113 0.021 ;
        RECT 5.223 -0.021 5.265 0.021 ;
        RECT 5.375 -0.021 5.417 0.021 ;
        RECT 0.435 0.149 0.477 0.191 ;
        RECT 0.739 0.149 0.781 0.191 ;
        RECT 1.043 0.149 1.085 0.191 ;
        RECT 1.347 0.149 1.389 0.191 ;
        RECT 1.651 0.149 1.693 0.191 ;
        RECT 1.955 0.149 1.997 0.191 ;
        RECT 2.259 0.149 2.301 0.191 ;
        RECT 2.563 0.149 2.605 0.191 ;
        RECT 2.867 0.149 2.909 0.191 ;
        RECT 3.171 0.149 3.213 0.191 ;
        RECT 3.475 0.149 3.517 0.191 ;
        RECT 3.779 0.149 3.821 0.191 ;
        RECT 4.083 0.149 4.125 0.191 ;
        RECT 4.387 0.149 4.429 0.191 ;
        RECT 4.691 0.149 4.733 0.191 ;
        RECT 4.995 0.149 5.037 0.191 ;
        RECT 0.435 0.241 0.477 0.283 ;
        RECT 0.739 0.241 0.781 0.283 ;
        RECT 1.043 0.241 1.085 0.283 ;
        RECT 1.347 0.241 1.389 0.283 ;
        RECT 1.651 0.241 1.693 0.283 ;
        RECT 1.955 0.241 1.997 0.283 ;
        RECT 2.259 0.241 2.301 0.283 ;
        RECT 2.563 0.241 2.605 0.283 ;
        RECT 2.867 0.241 2.909 0.283 ;
        RECT 3.171 0.241 3.213 0.283 ;
        RECT 3.475 0.241 3.517 0.283 ;
        RECT 3.779 0.241 3.821 0.283 ;
        RECT 4.083 0.241 4.125 0.283 ;
        RECT 4.387 0.241 4.429 0.283 ;
        RECT 4.691 0.241 4.733 0.283 ;
        RECT 4.995 0.241 5.037 0.283 ;
        RECT 0.435 0.333 0.477 0.375 ;
        RECT 0.739 0.333 0.781 0.375 ;
        RECT 1.043 0.333 1.085 0.375 ;
        RECT 1.347 0.333 1.389 0.375 ;
        RECT 1.651 0.333 1.693 0.375 ;
        RECT 1.955 0.333 1.997 0.375 ;
        RECT 2.259 0.333 2.301 0.375 ;
        RECT 2.563 0.333 2.605 0.375 ;
        RECT 2.867 0.333 2.909 0.375 ;
        RECT 3.171 0.333 3.213 0.375 ;
        RECT 3.475 0.333 3.517 0.375 ;
        RECT 3.779 0.333 3.821 0.375 ;
        RECT 4.083 0.333 4.125 0.375 ;
        RECT 4.387 0.333 4.429 0.375 ;
        RECT 4.691 0.333 4.733 0.375 ;
        RECT 4.995 0.333 5.037 0.375 ;
      LAYER M1 ;
        RECT 0 -0.03 5.472 0.03 ;
        RECT 2.863 0.03 2.913 0.41 ;
        RECT 3.167 0.03 3.217 0.41 ;
        RECT 3.471 0.03 3.521 0.41 ;
        RECT 3.775 0.03 3.825 0.41 ;
        RECT 4.079 0.03 4.129 0.41 ;
        RECT 4.383 0.03 4.433 0.41 ;
        RECT 4.687 0.03 4.737 0.41 ;
        RECT 4.991 0.03 5.041 0.41 ;
        RECT 0.431 0.03 0.481 0.41 ;
        RECT 0.735 0.03 0.785 0.41 ;
        RECT 1.039 0.03 1.089 0.41 ;
        RECT 1.343 0.03 1.393 0.41 ;
        RECT 1.647 0.03 1.697 0.41 ;
        RECT 1.951 0.03 2.001 0.41 ;
        RECT 2.255 0.03 2.305 0.41 ;
        RECT 2.559 0.03 2.609 0.41 ;
    END
  END VSS
  OBS
    LAYER PO ;
      RECT 5.381 0.069 5.411 1.606 ;
      RECT 5.229 0.069 5.259 1.606 ;
      RECT 5.077 0.069 5.107 1.606 ;
      RECT 4.925 0.069 4.955 1.606 ;
      RECT 4.621 0.069 4.651 1.606 ;
      RECT 4.773 0.069 4.803 1.606 ;
      RECT 4.317 0.069 4.347 1.606 ;
      RECT 4.469 0.069 4.499 1.606 ;
      RECT 4.165 0.069 4.195 1.606 ;
      RECT 4.013 0.069 4.043 1.606 ;
      RECT 3.861 0.069 3.891 1.606 ;
      RECT 3.709 0.069 3.739 1.606 ;
      RECT 3.405 0.069 3.435 1.606 ;
      RECT 3.557 0.069 3.587 1.606 ;
      RECT 2.797 0.069 2.827 1.606 ;
      RECT 2.949 0.069 2.979 1.606 ;
      RECT 2.645 0.069 2.675 1.606 ;
      RECT 3.101 0.069 3.131 1.606 ;
      RECT 3.253 0.069 3.283 1.606 ;
      RECT 1.429 0.069 1.459 1.606 ;
      RECT 1.581 0.069 1.611 1.606 ;
      RECT 1.733 0.069 1.763 1.606 ;
      RECT 2.341 0.069 2.371 1.606 ;
      RECT 2.189 0.069 2.219 1.606 ;
      RECT 2.037 0.069 2.067 1.606 ;
      RECT 1.885 0.069 1.915 1.606 ;
      RECT 2.493 0.069 2.523 1.606 ;
      RECT 1.277 0.069 1.307 1.606 ;
      RECT 1.125 0.069 1.155 1.606 ;
      RECT 0.973 0.069 1.003 1.606 ;
      RECT 0.213 0.069 0.243 1.606 ;
      RECT 0.365 0.069 0.395 1.606 ;
      RECT 0.821 0.069 0.851 1.606 ;
      RECT 0.669 0.069 0.699 1.606 ;
      RECT 0.517 0.069 0.547 1.606 ;
      RECT 0.061 0.069 0.091 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 5.587 1.773 ;
  END
END INVX32_RVT

MACRO AOI22X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.744 0.401 0.786 ;
      LAYER M1 ;
        RECT 0.249 0.705 0.404 0.815 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.932 0.553 0.974 ;
      LAYER M1 ;
        RECT 0.401 1.009 0.557 1.119 ;
        RECT 0.507 0.912 0.557 1.009 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.135 0.857 0.177 ;
      LAYER M1 ;
        RECT 0.705 0.097 0.863 0.207 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.6 0.705 0.642 ;
      LAYER M1 ;
        RECT 0.553 0.553 0.708 0.663 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 ;
  END A4
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.499 0.155 1.541 0.197 ;
        RECT 1.499 0.247 1.541 0.289 ;
        RECT 1.499 0.339 1.541 0.381 ;
        RECT 1.499 0.431 1.541 0.473 ;
        RECT 1.499 0.859 1.541 0.901 ;
        RECT 1.499 0.951 1.541 0.993 ;
        RECT 1.499 1.043 1.541 1.085 ;
        RECT 1.499 1.135 1.541 1.177 ;
        RECT 1.499 1.227 1.541 1.269 ;
        RECT 1.499 1.319 1.541 1.361 ;
        RECT 1.499 1.411 1.541 1.453 ;
      LAYER M1 ;
        RECT 1.495 1.271 1.545 1.473 ;
        RECT 1.465 1.161 1.575 1.271 ;
        RECT 1.495 0.854 1.545 1.161 ;
        RECT 1.495 0.804 1.585 0.854 ;
        RECT 1.535 0.493 1.585 0.804 ;
        RECT 1.495 0.443 1.585 0.493 ;
        RECT 1.495 0.135 1.545 0.443 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.043 1.134 1.085 1.176 ;
        RECT 1.347 1.217 1.389 1.259 ;
        RECT 1.043 1.226 1.085 1.268 ;
        RECT 1.347 1.309 1.389 1.351 ;
        RECT 1.043 1.318 1.085 1.36 ;
        RECT 1.347 1.401 1.389 1.443 ;
        RECT 0.435 1.407 0.477 1.449 ;
        RECT 1.043 1.41 1.085 1.452 ;
        RECT 1.347 1.493 1.389 1.535 ;
        RECT 0.435 1.499 0.477 1.541 ;
        RECT 1.043 1.502 1.085 1.544 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.824 1.702 ;
        RECT 0.431 1.387 0.481 1.642 ;
        RECT 1.039 1.114 1.089 1.642 ;
        RECT 1.342 1.197 1.392 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.347 0.135 1.389 0.177 ;
        RECT 1.347 0.227 1.389 0.269 ;
        RECT 0.587 0.315 0.629 0.357 ;
        RECT 1.347 0.319 1.389 0.361 ;
        RECT 1.043 0.409 1.085 0.451 ;
        RECT 1.347 0.411 1.389 0.453 ;
        RECT 1.043 0.501 1.085 0.543 ;
      LAYER M1 ;
        RECT 1.039 0.03 1.089 0.563 ;
        RECT 1.343 0.03 1.393 0.473 ;
        RECT 0.583 0.03 0.633 0.377 ;
        RECT 0 -0.03 1.824 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.191 0.612 1.485 0.662 ;
      RECT 1.191 1.003 1.396 1.053 ;
      RECT 1.346 0.662 1.396 1.003 ;
      RECT 1.191 1.053 1.241 1.564 ;
      RECT 1.191 1.002 1.241 1.003 ;
      RECT 1.191 0.662 1.241 0.663 ;
      RECT 1.191 0.389 1.241 0.612 ;
      RECT 0.887 1.337 0.937 1.571 ;
      RECT 0.583 1.337 0.633 1.571 ;
      RECT 0.279 1.287 0.937 1.337 ;
      RECT 0.279 1.337 0.329 1.571 ;
      RECT 0.735 0.846 1.181 0.896 ;
      RECT 0.279 0.279 0.329 0.452 ;
      RECT 0.887 0.279 0.937 0.452 ;
      RECT 0.279 0.452 0.937 0.502 ;
      RECT 0.758 0.502 0.808 0.813 ;
      RECT 0.735 0.813 0.808 0.846 ;
      RECT 0.735 0.896 0.785 1.237 ;
    LAYER PO ;
      RECT 1.581 0.064 1.611 1.605 ;
      RECT 1.429 0.065 1.459 1.605 ;
      RECT 0.213 0.072 0.243 1.621 ;
      RECT 0.821 0.072 0.851 1.621 ;
      RECT 1.733 0.064 1.763 1.605 ;
      RECT 0.973 0.076 1.003 1.621 ;
      RECT 1.277 0.06 1.307 1.614 ;
      RECT 0.061 0.072 0.091 1.621 ;
      RECT 0.365 0.067 0.395 1.621 ;
      RECT 0.517 0.072 0.547 1.621 ;
      RECT 0.669 0.072 0.699 1.621 ;
      RECT 1.125 0.06 1.155 1.614 ;
    LAYER CO ;
      RECT 0.891 0.299 0.933 0.341 ;
      RECT 0.587 1.325 0.629 1.367 ;
      RECT 0.587 1.417 0.629 1.459 ;
      RECT 0.739 1.083 0.781 1.125 ;
      RECT 0.739 1.175 0.781 1.217 ;
      RECT 0.283 1.417 0.325 1.459 ;
      RECT 0.283 1.325 0.325 1.367 ;
      RECT 0.283 1.509 0.325 1.551 ;
      RECT 0.283 0.299 0.325 0.341 ;
      RECT 1.195 0.409 1.237 0.451 ;
      RECT 0.587 1.509 0.629 1.551 ;
      RECT 1.423 0.616 1.465 0.658 ;
      RECT 1.119 0.85 1.161 0.892 ;
      RECT 1.195 0.501 1.237 0.543 ;
      RECT 1.195 1.502 1.237 1.544 ;
      RECT 0.891 1.325 0.933 1.367 ;
      RECT 0.891 1.509 0.933 1.551 ;
      RECT 1.195 1.318 1.237 1.36 ;
      RECT 1.195 1.226 1.237 1.268 ;
      RECT 0.283 0.391 0.325 0.433 ;
      RECT 1.195 1.41 1.237 1.452 ;
      RECT 0.891 0.391 0.933 0.433 ;
      RECT 1.195 1.134 1.237 1.176 ;
      RECT 0.891 1.417 0.933 1.459 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.939 1.773 ;
  END
END AOI22X1_RVT

MACRO OA21X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.271 0.81 0.421 0.817 ;
        RECT 0.249 0.717 0.421 0.81 ;
        RECT 0.249 0.701 0.359 0.717 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.027 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.482 0.553 1.524 ;
      LAYER M1 ;
        RECT 0.4 1.571 0.512 1.577 ;
        RECT 0.4 1.461 0.573 1.571 ;
        RECT 0.426 1.46 0.573 1.461 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.027 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.827 0.857 0.869 ;
      LAYER M1 ;
        RECT 0.712 0.962 0.861 0.986 ;
        RECT 0.705 0.853 0.861 0.962 ;
        RECT 0.811 0.807 0.861 0.853 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0135 ;
  END A3
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.195 0.239 1.237 0.281 ;
        RECT 1.195 0.331 1.237 0.373 ;
        RECT 1.195 0.423 1.237 0.465 ;
        RECT 1.195 0.987 1.237 1.029 ;
        RECT 1.195 1.079 1.237 1.121 ;
        RECT 1.195 1.171 1.237 1.213 ;
        RECT 1.195 1.263 1.237 1.305 ;
        RECT 1.195 1.355 1.237 1.397 ;
      LAYER M1 ;
        RECT 1.191 1.006 1.241 1.426 ;
        RECT 1.191 0.956 1.38 1.006 ;
        RECT 1.33 0.542 1.38 0.956 ;
        RECT 1.191 0.53 1.38 0.542 ;
        RECT 1.191 0.492 1.439 0.53 ;
        RECT 1.191 0.188 1.241 0.492 ;
        RECT 1.303 0.392 1.439 0.492 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 0.987 0.325 1.029 ;
        RECT 0.283 1.079 0.325 1.121 ;
        RECT 0.283 1.171 0.325 1.213 ;
        RECT 1.043 1.171 1.085 1.213 ;
        RECT 0.283 1.263 0.325 1.305 ;
        RECT 0.891 1.263 0.933 1.305 ;
        RECT 1.043 1.263 1.085 1.305 ;
        RECT 0.283 1.355 0.325 1.397 ;
        RECT 0.891 1.355 0.933 1.397 ;
        RECT 1.043 1.355 1.085 1.397 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.52 1.702 ;
        RECT 0.279 0.958 0.329 1.642 ;
        RECT 0.887 1.243 0.937 1.642 ;
        RECT 1.039 1.133 1.089 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.043 0.203 1.085 0.245 ;
        RECT 0.435 0.239 0.477 0.281 ;
        RECT 1.043 0.295 1.085 0.337 ;
        RECT 0.435 0.331 0.477 0.373 ;
        RECT 0.435 0.423 0.477 0.465 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.512 ;
        RECT 1.039 0.03 1.089 0.399 ;
        RECT 0 -0.03 1.52 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.079 0.681 1.165 0.699 ;
      RECT 1.079 0.613 1.165 0.631 ;
      RECT 0.887 0.631 1.176 0.681 ;
      RECT 0.583 1.18 0.633 1.393 ;
      RECT 0.583 1.106 0.633 1.13 ;
      RECT 0.735 1.18 0.785 1.393 ;
      RECT 0.735 1.106 0.785 1.13 ;
      RECT 0.913 0.681 0.963 1.13 ;
      RECT 0.887 0.181 0.937 0.631 ;
      RECT 0.583 1.13 0.963 1.18 ;
      RECT 0.279 0.598 0.633 0.648 ;
      RECT 0.735 0.181 0.785 0.412 ;
      RECT 0.583 0.412 0.785 0.462 ;
      RECT 0.583 0.462 0.633 0.598 ;
      RECT 0.583 0.181 0.633 0.412 ;
      RECT 0.279 0.178 0.329 0.598 ;
    LAYER PO ;
      RECT 0.973 0.101 1.003 1.469 ;
      RECT 0.365 0.101 0.395 1.469 ;
      RECT 0.821 0.101 0.851 1.469 ;
      RECT 1.277 0.101 1.307 1.469 ;
      RECT 1.429 0.101 1.459 1.469 ;
      RECT 0.061 0.101 0.091 1.469 ;
      RECT 1.125 0.069 1.155 1.608 ;
      RECT 0.517 0.101 0.547 1.567 ;
      RECT 0.213 0.101 0.243 1.469 ;
      RECT 0.669 0.101 0.699 1.469 ;
    LAYER CO ;
      RECT 0.283 0.239 0.325 0.281 ;
      RECT 0.739 1.23 0.781 1.272 ;
      RECT 0.739 1.322 0.781 1.364 ;
      RECT 0.587 0.423 0.629 0.465 ;
      RECT 0.283 0.423 0.325 0.465 ;
      RECT 0.283 0.331 0.325 0.373 ;
      RECT 0.739 0.303 0.781 0.345 ;
      RECT 0.739 0.211 0.781 0.253 ;
      RECT 0.587 1.23 0.629 1.272 ;
      RECT 0.587 1.322 0.629 1.364 ;
      RECT 0.587 1.138 0.629 1.18 ;
      RECT 0.587 0.239 0.629 0.281 ;
      RECT 0.587 0.331 0.629 0.373 ;
      RECT 1.119 0.635 1.161 0.677 ;
      RECT 0.891 0.211 0.933 0.253 ;
      RECT 0.891 0.303 0.933 0.345 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.635 1.787 ;
  END
END OA21X1_RVT

MACRO OAI221X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.271 0.81 0.421 0.817 ;
        RECT 0.249 0.71 0.421 0.81 ;
        RECT 0.249 0.701 0.359 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0222 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.482 0.553 1.524 ;
      LAYER M1 ;
        RECT 0.401 1.571 0.511 1.575 ;
        RECT 0.401 1.461 0.573 1.571 ;
        RECT 0.426 1.46 0.573 1.461 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0222 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.866 0.857 0.908 ;
      LAYER M1 ;
        RECT 0.811 1.002 0.968 1.139 ;
        RECT 0.811 0.842 0.861 1.002 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0222 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.739 0.705 0.781 ;
      LAYER M1 ;
        RECT 0.56 0.963 0.709 0.986 ;
        RECT 0.553 0.854 0.709 0.963 ;
        RECT 0.659 0.713 0.709 0.854 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0222 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.119 0.739 1.161 0.781 ;
      LAYER M1 ;
        RECT 1.115 0.675 1.165 0.808 ;
        RECT 1.023 0.658 1.165 0.675 ;
        RECT 1.009 0.601 1.165 0.658 ;
        RECT 1.009 0.549 1.123 0.601 ;
        RECT 1.023 0.541 1.123 0.549 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0162 ;
  END A5
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.803 0.239 1.845 0.281 ;
        RECT 1.803 0.331 1.845 0.373 ;
        RECT 1.803 0.423 1.845 0.465 ;
        RECT 1.803 0.987 1.845 1.029 ;
        RECT 1.803 1.079 1.845 1.121 ;
        RECT 1.803 1.171 1.845 1.213 ;
        RECT 1.803 1.263 1.845 1.305 ;
        RECT 1.803 1.355 1.845 1.397 ;
      LAYER M1 ;
        RECT 1.799 1.006 1.849 1.426 ;
        RECT 1.799 0.956 1.988 1.006 ;
        RECT 1.938 0.542 1.988 0.956 ;
        RECT 1.799 0.53 1.988 0.542 ;
        RECT 1.799 0.492 2.063 0.53 ;
        RECT 1.799 0.188 1.849 0.492 ;
        RECT 1.903 0.392 2.063 0.492 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.079 0.325 1.121 ;
        RECT 0.283 1.171 0.325 1.213 ;
        RECT 1.651 1.171 1.693 1.213 ;
        RECT 0.283 1.263 0.325 1.305 ;
        RECT 1.347 1.263 1.389 1.305 ;
        RECT 1.651 1.263 1.693 1.305 ;
        RECT 0.283 1.355 0.325 1.397 ;
        RECT 0.891 1.355 0.933 1.397 ;
        RECT 1.043 1.355 1.085 1.397 ;
        RECT 1.347 1.355 1.389 1.397 ;
        RECT 1.651 1.355 1.693 1.397 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 2.128 1.702 ;
        RECT 0.279 0.958 0.329 1.642 ;
        RECT 0.887 1.335 0.937 1.642 ;
        RECT 1.039 1.333 1.089 1.642 ;
        RECT 1.343 1.234 1.393 1.642 ;
        RECT 1.647 1.133 1.697 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 1.347 0.186 1.389 0.228 ;
        RECT 1.651 0.203 1.693 0.245 ;
        RECT 0.435 0.239 0.477 0.281 ;
        RECT 1.347 0.278 1.389 0.32 ;
        RECT 1.651 0.295 1.693 0.337 ;
        RECT 0.435 0.331 0.477 0.373 ;
        RECT 1.347 0.37 1.389 0.412 ;
        RECT 0.435 0.423 0.477 0.465 ;
      LAYER M1 ;
        RECT 1.343 0.03 1.393 0.532 ;
        RECT 0.431 0.03 0.481 0.512 ;
        RECT 1.647 0.03 1.697 0.399 ;
        RECT 0 -0.03 2.128 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.687 0.681 1.773 0.699 ;
      RECT 1.687 0.613 1.773 0.631 ;
      RECT 1.535 0.631 1.773 0.681 ;
      RECT 1.535 0.681 1.585 0.956 ;
      RECT 1.535 0.542 1.585 0.631 ;
      RECT 1.495 0.956 1.585 1.006 ;
      RECT 1.495 1.006 1.545 1.426 ;
      RECT 1.495 0.188 1.545 0.492 ;
      RECT 1.495 0.492 1.585 0.542 ;
      RECT 1.039 0.903 1.432 0.953 ;
      RECT 1.382 0.803 1.432 0.903 ;
      RECT 1.382 0.717 1.469 0.803 ;
      RECT 0.583 1.263 0.633 1.393 ;
      RECT 0.583 1.106 0.633 1.213 ;
      RECT 1.191 0.483 1.277 0.533 ;
      RECT 1.191 0.953 1.241 1.427 ;
      RECT 1.227 0.533 1.277 0.903 ;
      RECT 1.191 0.211 1.241 0.483 ;
      RECT 1.039 0.953 1.089 1.213 ;
      RECT 0.583 1.213 1.089 1.263 ;
      RECT 0.279 0.598 0.937 0.648 ;
      RECT 0.887 0.208 0.937 0.598 ;
      RECT 0.583 0.181 0.633 0.598 ;
      RECT 0.279 0.178 0.329 0.598 ;
      RECT 0.735 0.098 1.089 0.148 ;
      RECT 1.039 0.148 1.089 0.431 ;
      RECT 0.735 0.148 0.785 0.501 ;
    LAYER PO ;
      RECT 0.973 0.101 1.003 1.469 ;
      RECT 0.061 0.101 0.091 1.469 ;
      RECT 2.037 0.101 2.067 1.469 ;
      RECT 1.885 0.101 1.915 1.469 ;
      RECT 1.277 0.101 1.307 1.469 ;
      RECT 0.365 0.101 0.395 1.469 ;
      RECT 1.581 0.101 1.611 1.469 ;
      RECT 1.125 0.101 1.155 1.469 ;
      RECT 1.733 0.069 1.763 1.608 ;
      RECT 0.213 0.101 0.243 1.469 ;
      RECT 0.517 0.101 0.547 1.567 ;
      RECT 1.429 0.054 1.459 1.608 ;
      RECT 0.669 0.101 0.699 1.469 ;
      RECT 0.821 0.101 0.851 1.469 ;
    LAYER CO ;
      RECT 1.727 0.635 1.769 0.677 ;
      RECT 0.587 0.423 0.629 0.465 ;
      RECT 1.195 0.362 1.237 0.404 ;
      RECT 1.499 1.079 1.541 1.121 ;
      RECT 0.739 0.239 0.781 0.281 ;
      RECT 1.499 1.171 1.541 1.213 ;
      RECT 0.283 0.331 0.325 0.373 ;
      RECT 1.043 0.362 1.085 0.404 ;
      RECT 0.587 1.322 0.629 1.364 ;
      RECT 1.499 0.239 1.541 0.281 ;
      RECT 1.499 1.263 1.541 1.305 ;
      RECT 1.195 0.27 1.237 0.312 ;
      RECT 0.891 0.331 0.933 0.373 ;
      RECT 0.283 0.423 0.325 0.465 ;
      RECT 1.043 0.178 1.085 0.22 ;
      RECT 1.043 0.27 1.085 0.312 ;
      RECT 0.891 0.239 0.933 0.281 ;
      RECT 0.891 0.423 0.933 0.465 ;
      RECT 1.499 0.331 1.541 0.373 ;
      RECT 1.195 1.263 1.237 1.305 ;
      RECT 1.195 1.355 1.237 1.397 ;
      RECT 0.587 0.331 0.629 0.373 ;
      RECT 0.739 0.331 0.781 0.373 ;
      RECT 0.587 1.23 0.629 1.272 ;
      RECT 1.499 1.355 1.541 1.397 ;
      RECT 0.587 1.138 0.629 1.18 ;
      RECT 1.423 0.739 1.465 0.781 ;
      RECT 0.739 0.423 0.781 0.465 ;
      RECT 0.283 0.239 0.325 0.281 ;
      RECT 0.587 0.239 0.629 0.281 ;
    LAYER NWELL ;
      RECT -0.135 0.679 2.244 1.787 ;
  END
END OAI221X1_RVT

MACRO AO222X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.859 0.401 0.901 ;
      LAYER M1 ;
        RECT 0.247 0.857 0.421 0.967 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0249 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.6 0.553 0.642 ;
      LAYER M1 ;
        RECT 0.399 0.553 0.556 0.663 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0249 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.136 0.857 0.178 ;
      LAYER M1 ;
        RECT 0.703 0.097 0.863 0.207 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0249 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.857 0.705 0.899 ;
      LAYER M1 ;
        RECT 0.551 1.112 0.661 1.119 ;
        RECT 0.551 1.009 0.662 1.112 ;
        RECT 0.612 0.903 0.662 1.009 ;
        RECT 0.612 0.853 0.725 0.903 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0249 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.119 0.777 1.161 0.819 ;
      LAYER M1 ;
        RECT 1.007 0.773 1.181 0.823 ;
        RECT 1.007 0.705 1.117 0.773 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0249 ;
  END A5
  PIN A6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.271 0.543 1.313 0.585 ;
      LAYER M1 ;
        RECT 1.159 0.539 1.333 0.589 ;
        RECT 1.159 0.359 1.209 0.539 ;
        RECT 1.159 0.249 1.269 0.359 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0249 ;
  END A6
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.651 0.146 1.693 0.188 ;
        RECT 1.651 0.238 1.693 0.28 ;
        RECT 1.651 0.33 1.693 0.372 ;
        RECT 1.651 0.422 1.693 0.464 ;
        RECT 1.651 0.86 1.693 0.902 ;
        RECT 1.651 0.952 1.693 0.994 ;
        RECT 1.651 1.044 1.693 1.086 ;
        RECT 1.651 1.136 1.693 1.178 ;
        RECT 1.651 1.228 1.693 1.27 ;
        RECT 1.651 1.32 1.693 1.362 ;
        RECT 1.651 1.412 1.693 1.454 ;
        RECT 1.651 1.504 1.693 1.546 ;
      LAYER M1 ;
        RECT 1.647 1.271 1.697 1.566 ;
        RECT 1.615 1.161 1.725 1.271 ;
        RECT 1.647 0.865 1.697 1.161 ;
        RECT 1.647 0.864 1.737 0.865 ;
        RECT 1.647 0.815 1.747 0.864 ;
        RECT 1.697 0.484 1.747 0.815 ;
        RECT 1.647 0.434 1.747 0.484 ;
        RECT 1.647 0.126 1.697 0.434 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.499 1.044 1.541 1.086 ;
        RECT 1.499 1.136 1.541 1.178 ;
        RECT 1.499 1.228 1.541 1.27 ;
        RECT 1.499 1.32 1.541 1.362 ;
        RECT 0.435 1.407 0.477 1.449 ;
        RECT 1.499 1.412 1.541 1.454 ;
        RECT 0.435 1.499 0.477 1.541 ;
        RECT 1.499 1.504 1.541 1.546 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.976 1.702 ;
        RECT 0.431 1.387 0.481 1.642 ;
        RECT 1.495 1.024 1.545 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 1.499 0.146 1.541 0.188 ;
        RECT 1.499 0.238 1.541 0.28 ;
        RECT 1.347 0.312 1.389 0.354 ;
        RECT 0.587 0.326 0.629 0.368 ;
        RECT 1.499 0.33 1.541 0.372 ;
        RECT 1.347 0.404 1.389 0.446 ;
        RECT 0.587 0.418 0.629 0.46 ;
        RECT 1.499 0.422 1.541 0.464 ;
      LAYER M1 ;
        RECT 1.495 0.03 1.545 0.484 ;
        RECT 0.583 0.03 0.633 0.48 ;
        RECT 1.343 0.03 1.393 0.466 ;
        RECT 0 -0.03 1.976 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.461 0.636 1.637 0.686 ;
      RECT 1.19 0.907 1.511 0.908 ;
      RECT 0.887 0.908 1.511 0.957 ;
      RECT 1.461 0.686 1.511 0.907 ;
      RECT 0.279 0.318 0.329 0.713 ;
      RECT 0.887 0.957 1.24 0.958 ;
      RECT 1.19 0.958 1.24 1.484 ;
      RECT 1.039 0.363 1.089 0.487 ;
      RECT 0.887 0.313 1.089 0.363 ;
      RECT 0.887 0.763 0.937 0.908 ;
      RECT 0.279 0.713 0.937 0.763 ;
      RECT 0.887 0.363 0.937 0.713 ;
      RECT 1.342 1.208 1.392 1.534 ;
      RECT 1.039 1.071 1.089 1.534 ;
      RECT 1.039 1.534 1.392 1.584 ;
      RECT 0.735 1.071 0.785 1.237 ;
      RECT 0.755 1.021 1.089 1.025 ;
      RECT 0.735 1.025 1.089 1.071 ;
      RECT 0.583 1.337 0.633 1.571 ;
      RECT 0.279 1.287 0.937 1.337 ;
      RECT 0.887 1.337 0.937 1.571 ;
      RECT 0.279 1.337 0.329 1.571 ;
    LAYER PO ;
      RECT 1.733 0.075 1.763 1.616 ;
      RECT 1.429 0.075 1.459 1.616 ;
      RECT 1.277 0.076 1.307 1.621 ;
      RECT 0.669 0.072 0.699 1.621 ;
      RECT 0.517 0.072 0.547 1.621 ;
      RECT 0.365 0.067 0.395 1.621 ;
      RECT 1.885 0.075 1.915 1.616 ;
      RECT 0.061 0.072 0.091 1.621 ;
      RECT 0.973 0.076 1.003 1.621 ;
      RECT 1.581 0.076 1.611 1.616 ;
      RECT 0.821 0.072 0.851 1.621 ;
      RECT 0.213 0.072 0.243 1.621 ;
      RECT 1.125 0.076 1.155 1.621 ;
    LAYER CO ;
      RECT 0.587 1.417 0.629 1.459 ;
      RECT 0.587 1.325 0.629 1.367 ;
      RECT 0.283 0.43 0.325 0.472 ;
      RECT 0.891 0.428 0.933 0.47 ;
      RECT 0.891 1.509 0.933 1.551 ;
      RECT 1.575 0.639 1.617 0.681 ;
      RECT 0.891 0.336 0.933 0.378 ;
      RECT 0.283 0.338 0.325 0.38 ;
      RECT 0.891 1.417 0.933 1.459 ;
      RECT 1.195 1.238 1.237 1.28 ;
      RECT 1.195 1.33 1.237 1.372 ;
      RECT 1.195 1.146 1.237 1.188 ;
      RECT 1.195 1.422 1.237 1.464 ;
      RECT 1.043 1.504 1.085 1.546 ;
      RECT 1.043 0.425 1.085 0.467 ;
      RECT 1.043 0.333 1.085 0.375 ;
      RECT 1.043 1.32 1.085 1.362 ;
      RECT 1.043 1.412 1.085 1.454 ;
      RECT 0.283 1.325 0.325 1.367 ;
      RECT 1.347 1.228 1.389 1.27 ;
      RECT 1.347 1.32 1.389 1.362 ;
      RECT 1.347 1.412 1.389 1.454 ;
      RECT 1.347 1.504 1.389 1.546 ;
      RECT 1.043 1.228 1.085 1.27 ;
      RECT 1.043 1.136 1.085 1.178 ;
      RECT 0.891 1.325 0.933 1.367 ;
      RECT 0.587 1.509 0.629 1.551 ;
      RECT 0.283 1.417 0.325 1.459 ;
      RECT 0.283 1.509 0.325 1.551 ;
      RECT 0.739 1.175 0.781 1.217 ;
      RECT 0.739 1.083 0.781 1.125 ;
    LAYER NWELL ;
      RECT -0.115 0.679 2.091 1.773 ;
  END
END AO222X1_RVT

MACRO OA222X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.271 0.81 0.421 0.817 ;
        RECT 0.249 0.71 0.421 0.81 ;
        RECT 0.249 0.701 0.359 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.482 0.553 1.524 ;
      LAYER M1 ;
        RECT 0.401 1.571 0.511 1.575 ;
        RECT 0.401 1.461 0.573 1.571 ;
        RECT 0.426 1.46 0.573 1.461 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.866 0.857 0.908 ;
      LAYER M1 ;
        RECT 0.811 1.002 0.968 1.139 ;
        RECT 0.811 0.842 0.861 1.002 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.739 0.705 0.781 ;
      LAYER M1 ;
        RECT 0.56 0.963 0.709 0.986 ;
        RECT 0.553 0.854 0.709 0.963 ;
        RECT 0.659 0.713 0.709 0.854 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.119 0.739 1.161 0.781 ;
      LAYER M1 ;
        RECT 1.115 0.675 1.165 0.808 ;
        RECT 1.023 0.658 1.165 0.675 ;
        RECT 1.009 0.601 1.165 0.658 ;
        RECT 1.009 0.549 1.123 0.601 ;
        RECT 1.023 0.541 1.123 0.549 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A5
  PIN A6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.271 1.49 1.313 1.532 ;
      LAYER M1 ;
        RECT 1.171 1.485 1.339 1.535 ;
        RECT 1.171 1.281 1.221 1.485 ;
        RECT 1.171 1.266 1.28 1.281 ;
        RECT 1.16 1.157 1.28 1.266 ;
        RECT 1.171 1.146 1.28 1.157 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A6
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.651 0.239 1.693 0.281 ;
        RECT 1.651 0.331 1.693 0.373 ;
        RECT 1.651 0.423 1.693 0.465 ;
        RECT 1.651 0.987 1.693 1.029 ;
        RECT 1.651 1.079 1.693 1.121 ;
        RECT 1.651 1.171 1.693 1.213 ;
        RECT 1.651 1.263 1.693 1.305 ;
        RECT 1.651 1.355 1.693 1.397 ;
      LAYER M1 ;
        RECT 1.647 1.006 1.697 1.426 ;
        RECT 1.647 0.956 1.836 1.006 ;
        RECT 1.786 0.542 1.836 0.956 ;
        RECT 1.647 0.53 1.836 0.542 ;
        RECT 1.647 0.492 1.911 0.53 ;
        RECT 1.647 0.188 1.697 0.492 ;
        RECT 1.751 0.392 1.911 0.492 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.079 0.325 1.121 ;
        RECT 0.283 1.171 0.325 1.213 ;
        RECT 1.499 1.171 1.541 1.213 ;
        RECT 0.283 1.263 0.325 1.305 ;
        RECT 1.499 1.263 1.541 1.305 ;
        RECT 0.283 1.355 0.325 1.397 ;
        RECT 0.891 1.355 0.933 1.397 ;
        RECT 1.043 1.355 1.085 1.397 ;
        RECT 1.499 1.355 1.541 1.397 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.976 1.702 ;
        RECT 0.279 0.958 0.329 1.642 ;
        RECT 0.887 1.335 0.937 1.642 ;
        RECT 1.039 1.333 1.089 1.642 ;
        RECT 1.495 1.133 1.545 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 1.499 0.203 1.541 0.245 ;
        RECT 0.435 0.239 0.477 0.281 ;
        RECT 1.499 0.295 1.541 0.337 ;
        RECT 0.435 0.331 0.477 0.373 ;
        RECT 0.435 0.423 0.477 0.465 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.512 ;
        RECT 1.495 0.03 1.545 0.399 ;
        RECT 0 -0.03 1.976 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.343 0.631 1.621 0.681 ;
      RECT 1.535 0.681 1.621 0.699 ;
      RECT 1.535 0.613 1.621 0.631 ;
      RECT 0.583 1.263 0.633 1.393 ;
      RECT 0.583 1.106 0.633 1.213 ;
      RECT 1.039 0.903 1.393 0.953 ;
      RECT 1.191 0.483 1.393 0.533 ;
      RECT 1.343 0.533 1.393 0.631 ;
      RECT 1.343 0.953 1.393 1.38 ;
      RECT 1.343 0.681 1.393 0.903 ;
      RECT 1.191 0.211 1.241 0.483 ;
      RECT 1.039 0.953 1.089 1.213 ;
      RECT 0.583 1.213 1.089 1.263 ;
      RECT 0.279 0.598 0.937 0.648 ;
      RECT 0.887 0.208 0.937 0.598 ;
      RECT 0.583 0.181 0.633 0.598 ;
      RECT 0.279 0.178 0.329 0.598 ;
      RECT 1.343 0.148 1.393 0.432 ;
      RECT 0.735 0.098 1.393 0.148 ;
      RECT 1.039 0.148 1.089 0.431 ;
      RECT 0.735 0.148 0.785 0.501 ;
    LAYER PO ;
      RECT 1.277 0.101 1.307 1.567 ;
      RECT 1.581 0.069 1.611 1.608 ;
      RECT 1.125 0.101 1.155 1.469 ;
      RECT 1.429 0.101 1.459 1.469 ;
      RECT 0.365 0.101 0.395 1.469 ;
      RECT 1.885 0.101 1.915 1.469 ;
      RECT 0.061 0.101 0.091 1.469 ;
      RECT 1.733 0.101 1.763 1.469 ;
      RECT 0.973 0.101 1.003 1.469 ;
      RECT 0.821 0.101 0.851 1.469 ;
      RECT 0.669 0.101 0.699 1.469 ;
      RECT 0.517 0.101 0.547 1.567 ;
      RECT 0.213 0.101 0.243 1.469 ;
    LAYER CO ;
      RECT 1.195 0.362 1.237 0.404 ;
      RECT 0.283 0.331 0.325 0.373 ;
      RECT 0.283 0.239 0.325 0.281 ;
      RECT 1.575 0.635 1.617 0.677 ;
      RECT 0.739 0.331 0.781 0.373 ;
      RECT 0.587 1.138 0.629 1.18 ;
      RECT 0.587 1.322 0.629 1.364 ;
      RECT 0.587 1.23 0.629 1.272 ;
      RECT 0.587 0.331 0.629 0.373 ;
      RECT 1.347 0.178 1.389 0.22 ;
      RECT 0.587 0.239 0.629 0.281 ;
      RECT 1.347 0.27 1.389 0.312 ;
      RECT 1.043 0.178 1.085 0.22 ;
      RECT 1.043 0.27 1.085 0.312 ;
      RECT 1.347 1.289 1.389 1.331 ;
      RECT 1.347 1.197 1.389 1.239 ;
      RECT 0.283 0.423 0.325 0.465 ;
      RECT 0.587 0.423 0.629 0.465 ;
      RECT 1.195 0.27 1.237 0.312 ;
      RECT 0.739 0.423 0.781 0.465 ;
      RECT 1.347 0.362 1.389 0.404 ;
      RECT 0.891 0.423 0.933 0.465 ;
      RECT 0.891 0.331 0.933 0.373 ;
      RECT 0.891 0.239 0.933 0.281 ;
      RECT 1.043 0.362 1.085 0.404 ;
      RECT 0.739 0.239 0.781 0.281 ;
    LAYER NWELL ;
      RECT -0.135 0.679 2.092 1.787 ;
  END
END OA222X1_RVT

MACRO OA221X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.271 0.81 0.421 0.817 ;
        RECT 0.249 0.71 0.421 0.81 ;
        RECT 0.249 0.701 0.359 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0228 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.482 0.553 1.524 ;
      LAYER M1 ;
        RECT 0.401 1.571 0.511 1.577 ;
        RECT 0.401 1.461 0.573 1.571 ;
        RECT 0.426 1.46 0.573 1.461 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0228 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.866 0.857 0.908 ;
      LAYER M1 ;
        RECT 0.811 1.002 0.968 1.139 ;
        RECT 0.811 0.842 0.861 1.002 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0228 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.739 0.705 0.781 ;
      LAYER M1 ;
        RECT 0.56 0.963 0.709 0.986 ;
        RECT 0.553 0.854 0.709 0.963 ;
        RECT 0.659 0.713 0.709 0.854 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0228 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.119 0.739 1.161 0.781 ;
      LAYER M1 ;
        RECT 1.115 0.675 1.165 0.808 ;
        RECT 1.023 0.658 1.165 0.675 ;
        RECT 1.009 0.601 1.165 0.658 ;
        RECT 1.009 0.549 1.123 0.601 ;
        RECT 1.023 0.541 1.123 0.549 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0174 ;
  END A5
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.499 0.239 1.541 0.281 ;
        RECT 1.499 0.331 1.541 0.373 ;
        RECT 1.499 0.423 1.541 0.465 ;
        RECT 1.499 0.987 1.541 1.029 ;
        RECT 1.499 1.079 1.541 1.121 ;
        RECT 1.499 1.171 1.541 1.213 ;
        RECT 1.499 1.263 1.541 1.305 ;
        RECT 1.499 1.355 1.541 1.397 ;
      LAYER M1 ;
        RECT 1.495 1.006 1.545 1.426 ;
        RECT 1.495 0.956 1.684 1.006 ;
        RECT 1.634 0.542 1.684 0.956 ;
        RECT 1.495 0.53 1.684 0.542 ;
        RECT 1.495 0.492 1.759 0.53 ;
        RECT 1.495 0.188 1.545 0.492 ;
        RECT 1.599 0.392 1.759 0.492 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.079 0.325 1.121 ;
        RECT 0.283 1.171 0.325 1.213 ;
        RECT 1.347 1.171 1.389 1.213 ;
        RECT 0.283 1.263 0.325 1.305 ;
        RECT 1.347 1.263 1.389 1.305 ;
        RECT 0.283 1.355 0.325 1.397 ;
        RECT 0.891 1.355 0.933 1.397 ;
        RECT 1.043 1.355 1.085 1.397 ;
        RECT 1.347 1.355 1.389 1.397 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.824 1.702 ;
        RECT 0.279 0.958 0.329 1.642 ;
        RECT 0.887 1.335 0.937 1.642 ;
        RECT 1.039 1.333 1.089 1.642 ;
        RECT 1.343 1.133 1.393 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.347 0.203 1.389 0.245 ;
        RECT 0.435 0.239 0.477 0.281 ;
        RECT 1.347 0.295 1.389 0.337 ;
        RECT 0.435 0.331 0.477 0.373 ;
        RECT 0.435 0.423 0.477 0.465 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.512 ;
        RECT 1.343 0.03 1.393 0.399 ;
        RECT 0 -0.03 1.824 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.383 0.681 1.469 0.699 ;
      RECT 1.383 0.613 1.469 0.631 ;
      RECT 1.227 0.631 1.469 0.681 ;
      RECT 0.583 1.263 0.633 1.393 ;
      RECT 0.583 1.106 0.633 1.213 ;
      RECT 1.039 0.903 1.277 0.953 ;
      RECT 1.191 0.483 1.277 0.533 ;
      RECT 1.227 0.533 1.277 0.631 ;
      RECT 1.191 0.953 1.241 1.427 ;
      RECT 1.227 0.681 1.277 0.903 ;
      RECT 1.191 0.211 1.241 0.483 ;
      RECT 1.039 0.953 1.089 1.213 ;
      RECT 0.583 1.213 1.089 1.263 ;
      RECT 0.279 0.598 0.937 0.648 ;
      RECT 0.887 0.208 0.937 0.598 ;
      RECT 0.583 0.181 0.633 0.598 ;
      RECT 0.279 0.178 0.329 0.598 ;
      RECT 0.735 0.098 1.089 0.148 ;
      RECT 0.735 0.148 0.785 0.501 ;
      RECT 1.039 0.148 1.089 0.431 ;
    LAYER PO ;
      RECT 1.277 0.101 1.307 1.469 ;
      RECT 0.365 0.101 0.395 1.469 ;
      RECT 0.973 0.101 1.003 1.469 ;
      RECT 0.061 0.101 0.091 1.469 ;
      RECT 1.733 0.101 1.763 1.469 ;
      RECT 1.581 0.101 1.611 1.469 ;
      RECT 1.125 0.101 1.155 1.469 ;
      RECT 1.429 0.069 1.459 1.608 ;
      RECT 0.213 0.101 0.243 1.469 ;
      RECT 0.517 0.101 0.547 1.567 ;
      RECT 0.669 0.101 0.699 1.469 ;
      RECT 0.821 0.101 0.851 1.469 ;
    LAYER CO ;
      RECT 1.195 0.362 1.237 0.404 ;
      RECT 0.283 0.331 0.325 0.373 ;
      RECT 1.195 0.27 1.237 0.312 ;
      RECT 0.587 0.423 0.629 0.465 ;
      RECT 0.891 0.331 0.933 0.373 ;
      RECT 0.283 0.423 0.325 0.465 ;
      RECT 1.195 1.355 1.237 1.397 ;
      RECT 0.891 0.423 0.933 0.465 ;
      RECT 1.043 0.362 1.085 0.404 ;
      RECT 1.423 0.635 1.465 0.677 ;
      RECT 0.891 0.239 0.933 0.281 ;
      RECT 1.043 0.27 1.085 0.312 ;
      RECT 1.043 0.178 1.085 0.22 ;
      RECT 0.739 0.239 0.781 0.281 ;
      RECT 0.587 1.138 0.629 1.18 ;
      RECT 0.739 0.331 0.781 0.373 ;
      RECT 0.587 0.239 0.629 0.281 ;
      RECT 0.283 0.239 0.325 0.281 ;
      RECT 0.739 0.423 0.781 0.465 ;
      RECT 0.587 0.331 0.629 0.373 ;
      RECT 0.587 1.23 0.629 1.272 ;
      RECT 0.587 1.322 0.629 1.364 ;
      RECT 1.195 1.263 1.237 1.305 ;
    LAYER NWELL ;
      RECT -0.135 0.679 1.94 1.787 ;
  END
END OA221X1_RVT

MACRO NOR2X0_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.665 0.401 0.707 ;
      LAYER M1 ;
        RECT 0.249 0.631 0.421 0.815 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0303 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.665 0.553 0.707 ;
      LAYER M1 ;
        RECT 0.489 0.553 0.663 0.733 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0303 ;
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.195 0.151 1.237 0.193 ;
        RECT 1.195 0.245 1.237 0.287 ;
        RECT 1.195 0.337 1.237 0.379 ;
        RECT 1.195 0.43 1.237 0.472 ;
        RECT 1.195 0.841 1.237 0.883 ;
        RECT 1.195 0.933 1.237 0.975 ;
        RECT 1.195 1.027 1.237 1.069 ;
        RECT 1.195 1.119 1.237 1.161 ;
        RECT 1.195 1.212 1.237 1.254 ;
        RECT 1.195 1.304 1.237 1.346 ;
        RECT 1.195 1.398 1.237 1.44 ;
        RECT 1.195 1.49 1.237 1.532 ;
      LAYER M1 ;
        RECT 1.191 0.824 1.241 1.552 ;
        RECT 1.191 0.774 1.395 0.824 ;
        RECT 1.345 0.511 1.395 0.774 ;
        RECT 1.313 0.49 1.423 0.511 ;
        RECT 1.191 0.49 1.241 0.492 ;
        RECT 1.191 0.44 1.423 0.49 ;
        RECT 1.191 0.131 1.241 0.44 ;
        RECT 1.313 0.401 1.423 0.44 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 0.931 0.325 0.973 ;
        RECT 1.043 0.931 1.085 0.973 ;
        RECT 0.739 1.008 0.781 1.05 ;
        RECT 0.283 1.024 0.325 1.066 ;
        RECT 1.043 1.024 1.085 1.066 ;
        RECT 0.739 1.1 0.781 1.142 ;
        RECT 0.283 1.116 0.325 1.158 ;
        RECT 1.043 1.116 1.085 1.158 ;
        RECT 0.283 1.209 0.325 1.251 ;
        RECT 1.043 1.209 1.085 1.251 ;
        RECT 0.283 1.301 0.325 1.343 ;
        RECT 1.043 1.301 1.085 1.343 ;
        RECT 0.283 1.395 0.325 1.437 ;
        RECT 1.043 1.395 1.085 1.437 ;
        RECT 0.283 1.487 0.325 1.529 ;
        RECT 1.043 1.487 1.085 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.52 1.702 ;
        RECT 0.279 0.911 0.329 1.642 ;
        RECT 0.735 0.988 0.785 1.642 ;
        RECT 1.039 0.911 1.089 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 0.739 0.141 0.781 0.183 ;
        RECT 1.043 0.141 1.085 0.183 ;
        RECT 0.435 0.176 0.477 0.218 ;
        RECT 0.739 0.233 0.781 0.275 ;
        RECT 1.043 0.233 1.085 0.275 ;
        RECT 0.435 0.268 0.477 0.31 ;
        RECT 1.043 0.325 1.085 0.367 ;
      LAYER M1 ;
        RECT 1.039 0.03 1.089 0.387 ;
        RECT 0.431 0.03 0.481 0.33 ;
        RECT 0.735 0.03 0.785 0.295 ;
        RECT 0 -0.03 1.52 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.279 0.383 0.775 0.433 ;
      RECT 0.583 0.813 0.775 0.863 ;
      RECT 0.725 0.666 0.877 0.716 ;
      RECT 0.725 0.433 0.775 0.666 ;
      RECT 0.725 0.716 0.775 0.813 ;
      RECT 0.279 0.174 0.329 0.383 ;
      RECT 0.583 0.174 0.633 0.383 ;
      RECT 0.583 0.863 0.633 1.552 ;
      RECT 0.887 0.773 1.06 0.823 ;
      RECT 0.887 0.502 1.061 0.552 ;
      RECT 1.01 0.711 1.06 0.773 ;
      RECT 1.01 0.661 1.181 0.711 ;
      RECT 1.01 0.552 1.06 0.661 ;
      RECT 0.887 0.823 0.937 1.152 ;
      RECT 0.887 0.131 0.937 0.502 ;
    LAYER PO ;
      RECT 1.125 0.071 1.155 1.612 ;
      RECT 1.277 0.071 1.307 1.612 ;
      RECT 0.821 0.071 0.851 1.612 ;
      RECT 0.973 0.071 1.003 1.612 ;
      RECT 0.061 0.071 0.091 1.612 ;
      RECT 1.429 0.071 1.459 1.612 ;
      RECT 0.213 0.071 0.243 1.612 ;
      RECT 0.669 0.071 0.699 1.612 ;
      RECT 0.365 0.071 0.395 1.612 ;
      RECT 0.517 0.071 0.547 1.612 ;
    LAYER CO ;
      RECT 0.587 1.49 0.629 1.532 ;
      RECT 0.587 1.396 0.629 1.438 ;
      RECT 0.587 1.304 0.629 1.346 ;
      RECT 0.587 1.211 0.629 1.253 ;
      RECT 0.587 0.194 0.629 0.236 ;
      RECT 0.283 0.194 0.325 0.236 ;
      RECT 0.891 0.812 0.933 0.854 ;
      RECT 0.587 0.842 0.629 0.884 ;
      RECT 0.587 0.934 0.629 0.976 ;
      RECT 0.587 1.027 0.629 1.069 ;
      RECT 0.815 0.67 0.857 0.712 ;
      RECT 0.891 0.245 0.933 0.287 ;
      RECT 0.891 0.151 0.933 0.193 ;
      RECT 1.119 0.665 1.161 0.707 ;
      RECT 0.587 1.119 0.629 1.161 ;
      RECT 0.891 1.09 0.933 1.132 ;
      RECT 0.891 0.998 0.933 1.04 ;
      RECT 0.891 0.904 0.933 0.946 ;
      RECT 0.587 0.288 0.629 0.33 ;
      RECT 0.283 0.288 0.325 0.33 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.635 1.773 ;
  END
END NOR2X0_RVT

MACRO NAND2X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.891 0.553 0.933 ;
      LAYER M1 ;
        RECT 0.553 0.937 0.663 0.967 ;
        RECT 0.456 0.887 0.663 0.937 ;
        RECT 0.553 0.857 0.663 0.887 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.401 0.785 0.511 0.815 ;
        RECT 0.339 0.735 0.511 0.785 ;
        RECT 0.401 0.705 0.511 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.195 0.142 1.237 0.184 ;
        RECT 1.195 0.234 1.237 0.276 ;
        RECT 1.195 0.835 1.237 0.877 ;
        RECT 1.195 0.927 1.237 0.969 ;
        RECT 1.195 1.019 1.237 1.061 ;
        RECT 1.195 1.111 1.237 1.153 ;
        RECT 1.195 1.203 1.237 1.245 ;
        RECT 1.195 1.295 1.237 1.337 ;
        RECT 1.195 1.387 1.237 1.429 ;
        RECT 1.195 1.479 1.237 1.521 ;
      LAYER M1 ;
        RECT 1.191 0.792 1.241 1.556 ;
        RECT 1.191 0.742 1.515 0.792 ;
        RECT 1.465 0.663 1.515 0.742 ;
        RECT 1.465 0.592 1.575 0.663 ;
        RECT 1.191 0.553 1.575 0.592 ;
        RECT 1.191 0.542 1.515 0.553 ;
        RECT 1.191 0.114 1.241 0.542 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.043 0.835 1.085 0.877 ;
        RECT 1.043 0.927 1.085 0.969 ;
        RECT 1.347 0.927 1.389 0.969 ;
        RECT 1.043 1.019 1.085 1.061 ;
        RECT 1.347 1.019 1.389 1.061 ;
        RECT 1.043 1.111 1.085 1.153 ;
        RECT 1.347 1.111 1.389 1.153 ;
        RECT 0.739 1.203 0.781 1.245 ;
        RECT 1.043 1.203 1.085 1.245 ;
        RECT 1.347 1.203 1.389 1.245 ;
        RECT 0.435 1.213 0.477 1.255 ;
        RECT 0.739 1.295 0.781 1.337 ;
        RECT 1.043 1.295 1.085 1.337 ;
        RECT 1.347 1.295 1.389 1.337 ;
        RECT 0.435 1.305 0.477 1.347 ;
        RECT 0.739 1.387 0.781 1.429 ;
        RECT 1.043 1.387 1.085 1.429 ;
        RECT 1.347 1.387 1.389 1.429 ;
        RECT 0.435 1.397 0.477 1.439 ;
        RECT 0.739 1.479 0.781 1.521 ;
        RECT 1.043 1.479 1.085 1.521 ;
        RECT 1.347 1.479 1.389 1.521 ;
        RECT 0.435 1.489 0.477 1.531 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.672 1.702 ;
        RECT 0.431 1.193 0.481 1.642 ;
        RECT 0.735 1.183 0.785 1.642 ;
        RECT 1.039 0.815 1.089 1.642 ;
        RECT 1.343 0.907 1.393 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 0.283 0.141 0.325 0.183 ;
        RECT 0.739 0.142 0.781 0.184 ;
        RECT 1.043 0.142 1.085 0.184 ;
        RECT 1.347 0.142 1.389 0.184 ;
        RECT 0.283 0.233 0.325 0.275 ;
        RECT 0.739 0.234 0.781 0.276 ;
        RECT 1.043 0.234 1.085 0.276 ;
        RECT 1.347 0.234 1.389 0.276 ;
        RECT 0.283 0.325 0.325 0.367 ;
        RECT 1.043 0.326 1.085 0.368 ;
        RECT 1.347 0.326 1.389 0.368 ;
        RECT 0.283 0.417 0.325 0.459 ;
        RECT 1.043 0.418 1.085 0.46 ;
        RECT 1.347 0.418 1.389 0.46 ;
      LAYER M1 ;
        RECT 1.039 0.03 1.089 0.48 ;
        RECT 1.343 0.03 1.393 0.48 ;
        RECT 0.279 0.03 0.329 0.479 ;
        RECT 0.735 0.03 0.785 0.296 ;
        RECT 0 -0.03 1.672 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.587 0.141 0.629 0.183 ;
      RECT 0.587 0.233 0.629 0.275 ;
      RECT 1.271 0.646 1.313 0.688 ;
      RECT 0.587 0.325 0.629 0.367 ;
      RECT 0.587 0.417 0.629 0.459 ;
      RECT 0.891 0.142 0.933 0.184 ;
      RECT 0.891 1.203 0.933 1.245 ;
      RECT 0.815 0.735 0.857 0.777 ;
      RECT 1.119 0.646 1.161 0.688 ;
      RECT 0.891 0.142 0.933 0.184 ;
      RECT 0.891 1.479 0.933 1.521 ;
      RECT 0.891 0.234 0.933 0.276 ;
      RECT 0.891 1.387 0.933 1.429 ;
      RECT 0.891 1.295 0.933 1.337 ;
      RECT 0.891 1.203 0.933 1.245 ;
      RECT 0.891 1.479 0.933 1.521 ;
      RECT 0.587 1.489 0.629 1.531 ;
      RECT 0.587 1.397 0.629 1.439 ;
      RECT 0.587 1.305 0.629 1.347 ;
      RECT 0.587 1.213 0.629 1.255 ;
      RECT 0.283 1.213 0.325 1.255 ;
      RECT 0.283 1.305 0.325 1.347 ;
      RECT 0.283 1.489 0.325 1.531 ;
      RECT 0.283 1.397 0.325 1.439 ;
      RECT 0.891 1.387 0.933 1.429 ;
      RECT 0.891 1.295 0.933 1.337 ;
    LAYER M1 ;
      RECT 0.71 0.731 0.877 0.781 ;
      RECT 0.713 0.663 0.763 0.731 ;
      RECT 0.279 1.083 0.763 1.133 ;
      RECT 0.583 0.613 0.763 0.663 ;
      RECT 0.713 0.781 0.763 1.083 ;
      RECT 0.279 1.133 0.329 1.551 ;
      RECT 0.583 1.133 0.633 1.551 ;
      RECT 0.583 0.121 0.633 0.613 ;
      RECT 0.927 0.642 1.333 0.692 ;
      RECT 0.887 0.906 0.937 1.556 ;
      RECT 0.887 0.856 0.977 0.906 ;
      RECT 0.887 0.114 0.937 0.455 ;
      RECT 0.887 0.455 0.977 0.505 ;
      RECT 0.927 0.692 0.977 0.856 ;
      RECT 0.927 0.505 0.977 0.642 ;
    LAYER PO ;
      RECT 0.669 0.071 0.699 1.601 ;
      RECT 0.365 0.071 0.395 1.601 ;
      RECT 0.517 0.071 0.547 1.601 ;
      RECT 0.213 0.071 0.243 1.601 ;
      RECT 0.061 0.071 0.091 1.601 ;
      RECT 1.277 0.064 1.307 1.604 ;
      RECT 0.973 0.064 1.003 1.6 ;
      RECT 0.821 0.064 0.851 1.61 ;
      RECT 1.125 0.064 1.155 1.605 ;
      RECT 1.581 0.064 1.611 1.6 ;
      RECT 1.429 0.064 1.459 1.602 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.787 1.773 ;
  END
END NAND2X2_RVT

MACRO NAND3X4_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.739 0.705 0.781 ;
      LAYER M1 ;
        RECT 0.553 0.785 0.663 0.815 ;
        RECT 0.553 0.735 0.725 0.785 ;
        RECT 0.553 0.705 0.663 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.043 0.553 1.085 ;
      LAYER M1 ;
        RECT 0.401 1.089 0.511 1.119 ;
        RECT 0.401 1.039 0.573 1.089 ;
        RECT 0.401 1.009 0.511 1.039 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.737 0.401 0.779 ;
      LAYER M1 ;
        RECT 0.249 0.785 0.359 0.815 ;
        RECT 0.249 0.735 0.421 0.785 ;
        RECT 0.249 0.704 0.359 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END A3
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.195 0.15 1.237 0.192 ;
        RECT 1.499 0.15 1.541 0.192 ;
        RECT 1.803 0.152 1.845 0.194 ;
        RECT 1.195 0.242 1.237 0.284 ;
        RECT 1.499 0.242 1.541 0.284 ;
        RECT 1.803 0.244 1.845 0.286 ;
        RECT 1.195 0.334 1.237 0.376 ;
        RECT 1.499 0.334 1.541 0.376 ;
        RECT 1.803 0.336 1.845 0.378 ;
        RECT 1.195 0.426 1.237 0.468 ;
        RECT 1.499 0.426 1.541 0.468 ;
        RECT 1.803 0.428 1.845 0.47 ;
        RECT 1.195 0.844 1.237 0.886 ;
        RECT 1.499 0.844 1.541 0.886 ;
        RECT 1.803 0.844 1.845 0.886 ;
        RECT 1.195 0.936 1.237 0.978 ;
        RECT 1.499 0.936 1.541 0.978 ;
        RECT 1.803 0.936 1.845 0.978 ;
        RECT 1.195 1.028 1.237 1.07 ;
        RECT 1.499 1.028 1.541 1.07 ;
        RECT 1.803 1.028 1.845 1.07 ;
        RECT 1.195 1.12 1.237 1.162 ;
        RECT 1.499 1.12 1.541 1.162 ;
        RECT 1.803 1.12 1.845 1.162 ;
        RECT 1.195 1.212 1.237 1.254 ;
        RECT 1.499 1.212 1.541 1.254 ;
        RECT 1.803 1.212 1.845 1.254 ;
        RECT 1.195 1.304 1.237 1.346 ;
        RECT 1.499 1.304 1.541 1.346 ;
        RECT 1.803 1.304 1.845 1.346 ;
        RECT 1.195 1.396 1.237 1.438 ;
        RECT 1.499 1.396 1.541 1.438 ;
        RECT 1.803 1.396 1.845 1.438 ;
        RECT 1.195 1.488 1.237 1.53 ;
        RECT 1.499 1.488 1.541 1.53 ;
        RECT 1.803 1.488 1.845 1.53 ;
      LAYER M1 ;
        RECT 1.191 0.793 1.241 1.565 ;
        RECT 1.495 0.793 1.545 1.565 ;
        RECT 1.799 0.793 1.849 1.565 ;
        RECT 1.191 0.743 1.954 0.793 ;
        RECT 1.904 0.663 1.954 0.743 ;
        RECT 1.904 0.564 2.041 0.663 ;
        RECT 1.191 0.553 2.041 0.564 ;
        RECT 1.191 0.514 1.954 0.553 ;
        RECT 1.191 0.115 1.241 0.514 ;
        RECT 1.495 0.115 1.545 0.514 ;
        RECT 1.799 0.115 1.849 0.514 ;
    END
    ANTENNADIFFAREA 0.3972 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.347 0.936 1.389 0.978 ;
        RECT 1.651 0.936 1.693 0.978 ;
        RECT 1.347 1.028 1.389 1.07 ;
        RECT 1.651 1.028 1.693 1.07 ;
        RECT 1.347 1.12 1.389 1.162 ;
        RECT 1.651 1.12 1.693 1.162 ;
        RECT 0.891 1.203 0.933 1.245 ;
        RECT 1.347 1.212 1.389 1.254 ;
        RECT 1.651 1.212 1.693 1.254 ;
        RECT 0.891 1.295 0.933 1.337 ;
        RECT 1.347 1.304 1.389 1.346 ;
        RECT 1.651 1.304 1.693 1.346 ;
        RECT 0.891 1.387 0.933 1.429 ;
        RECT 1.347 1.396 1.389 1.438 ;
        RECT 1.651 1.396 1.693 1.438 ;
        RECT 0.283 1.397 0.325 1.439 ;
        RECT 0.587 1.397 0.629 1.439 ;
        RECT 0.891 1.479 0.933 1.521 ;
        RECT 1.347 1.488 1.389 1.53 ;
        RECT 1.651 1.488 1.693 1.53 ;
        RECT 0.283 1.489 0.325 1.531 ;
        RECT 0.587 1.489 0.629 1.531 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 2.128 1.702 ;
        RECT 0.279 1.377 0.329 1.642 ;
        RECT 0.583 1.377 0.633 1.642 ;
        RECT 0.887 1.183 0.937 1.642 ;
        RECT 1.343 0.847 1.393 1.642 ;
        RECT 1.647 0.847 1.697 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 0.283 0.141 0.325 0.183 ;
        RECT 0.891 0.142 0.933 0.184 ;
        RECT 1.347 0.152 1.389 0.194 ;
        RECT 1.651 0.152 1.693 0.194 ;
        RECT 0.283 0.233 0.325 0.275 ;
        RECT 0.891 0.234 0.933 0.276 ;
        RECT 1.347 0.244 1.389 0.286 ;
        RECT 1.651 0.244 1.693 0.286 ;
        RECT 0.283 0.325 0.325 0.367 ;
        RECT 1.347 0.336 1.389 0.378 ;
        RECT 1.651 0.336 1.693 0.378 ;
        RECT 0.283 0.417 0.325 0.459 ;
      LAYER M1 ;
        RECT 0.279 0.03 0.329 0.479 ;
        RECT 1.343 0.03 1.393 0.413 ;
        RECT 1.647 0.03 1.697 0.413 ;
        RECT 0.887 0.03 0.937 0.296 ;
        RECT 0 -0.03 2.128 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.435 1.489 0.477 1.531 ;
      RECT 0.739 1.489 0.781 1.531 ;
      RECT 0.739 0.325 0.781 0.367 ;
      RECT 1.043 1.387 1.085 1.429 ;
      RECT 1.043 1.387 1.085 1.429 ;
      RECT 1.043 1.203 1.085 1.245 ;
      RECT 1.043 1.295 1.085 1.337 ;
      RECT 1.043 1.479 1.085 1.521 ;
      RECT 1.043 1.203 1.085 1.245 ;
      RECT 0.739 1.397 0.781 1.439 ;
      RECT 0.739 0.417 0.781 0.459 ;
      RECT 0.435 1.397 0.477 1.439 ;
      RECT 0.739 0.233 0.781 0.275 ;
      RECT 0.739 0.141 0.781 0.183 ;
      RECT 1.043 1.295 1.085 1.337 ;
      RECT 0.967 0.735 1.009 0.777 ;
      RECT 1.575 0.646 1.617 0.688 ;
      RECT 1.271 0.646 1.313 0.688 ;
      RECT 1.727 0.646 1.769 0.688 ;
      RECT 1.423 0.646 1.465 0.688 ;
      RECT 1.043 0.234 1.085 0.276 ;
      RECT 1.043 0.142 1.085 0.184 ;
      RECT 1.043 0.142 1.085 0.184 ;
      RECT 1.043 1.479 1.085 1.521 ;
    LAYER M1 ;
      RECT 1.079 0.642 1.789 0.692 ;
      RECT 1.039 0.906 1.089 1.556 ;
      RECT 1.039 0.856 1.129 0.906 ;
      RECT 1.039 0.114 1.089 0.455 ;
      RECT 1.039 0.455 1.129 0.505 ;
      RECT 1.079 0.505 1.129 0.642 ;
      RECT 1.079 0.692 1.129 0.856 ;
      RECT 0.777 0.731 1.029 0.781 ;
      RECT 0.431 1.235 0.481 1.551 ;
      RECT 0.735 0.571 0.827 0.621 ;
      RECT 0.735 0.121 0.785 0.571 ;
      RECT 0.735 1.235 0.785 1.551 ;
      RECT 0.431 1.185 0.827 1.235 ;
      RECT 0.777 0.621 0.827 0.731 ;
      RECT 0.777 0.781 0.827 1.185 ;
    LAYER PO ;
      RECT 0.669 0.071 0.699 1.61 ;
      RECT 0.973 0.064 1.003 1.61 ;
      RECT 0.213 0.071 0.243 1.61 ;
      RECT 0.517 0.071 0.547 1.61 ;
      RECT 0.365 0.071 0.395 1.61 ;
      RECT 1.125 0.064 1.155 1.6 ;
      RECT 0.061 0.071 0.091 1.61 ;
      RECT 0.821 0.071 0.851 1.61 ;
      RECT 1.429 0.072 1.459 1.61 ;
      RECT 1.581 0.072 1.611 1.61 ;
      RECT 1.733 0.072 1.763 1.61 ;
      RECT 2.037 0.072 2.067 1.61 ;
      RECT 1.885 0.072 1.915 1.61 ;
      RECT 1.277 0.072 1.307 1.61 ;
    LAYER NWELL ;
      RECT -0.115 0.679 2.243 1.773 ;
  END
END NAND3X4_RVT

MACRO OR4X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.666 0.401 0.708 ;
      LAYER M1 ;
        RECT 0.249 0.662 0.421 0.712 ;
        RECT 0.249 0.553 0.359 0.662 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.666 0.553 0.708 ;
      LAYER M1 ;
        RECT 0.507 0.857 0.663 0.967 ;
        RECT 0.507 0.646 0.557 0.857 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.666 0.705 0.708 ;
      LAYER M1 ;
        RECT 0.659 0.511 0.709 0.728 ;
        RECT 0.659 0.401 0.815 0.511 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.666 0.857 0.708 ;
      LAYER M1 ;
        RECT 0.809 0.705 0.967 0.815 ;
        RECT 0.811 0.646 0.861 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A4
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.803 0.151 1.845 0.193 ;
        RECT 1.803 0.245 1.845 0.287 ;
        RECT 1.803 0.337 1.845 0.379 ;
        RECT 1.803 0.43 1.845 0.472 ;
        RECT 1.803 0.841 1.845 0.883 ;
        RECT 1.803 0.933 1.845 0.975 ;
        RECT 1.803 1.027 1.845 1.069 ;
        RECT 1.803 1.119 1.845 1.161 ;
        RECT 1.803 1.212 1.845 1.254 ;
        RECT 1.803 1.304 1.845 1.346 ;
        RECT 1.803 1.398 1.845 1.44 ;
        RECT 1.803 1.49 1.845 1.532 ;
      LAYER M1 ;
        RECT 1.799 0.838 1.849 1.552 ;
        RECT 1.799 0.788 2.159 0.838 ;
        RECT 2.109 0.553 2.159 0.788 ;
        RECT 1.799 0.503 2.159 0.553 ;
        RECT 1.799 0.131 1.849 0.503 ;
        RECT 2.109 0.359 2.159 0.503 ;
        RECT 2.073 0.249 2.183 0.359 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 0.838 0.325 0.88 ;
        RECT 0.283 0.93 0.325 0.972 ;
        RECT 1.955 0.931 1.997 0.973 ;
        RECT 1.347 0.932 1.389 0.974 ;
        RECT 1.651 0.932 1.693 0.974 ;
        RECT 0.283 1.024 0.325 1.066 ;
        RECT 1.347 1.024 1.389 1.066 ;
        RECT 1.651 1.024 1.693 1.066 ;
        RECT 1.955 1.024 1.997 1.066 ;
        RECT 1.043 1.085 1.085 1.127 ;
        RECT 0.283 1.116 0.325 1.158 ;
        RECT 1.347 1.116 1.389 1.158 ;
        RECT 1.651 1.116 1.693 1.158 ;
        RECT 1.955 1.116 1.997 1.158 ;
        RECT 0.283 1.209 0.325 1.251 ;
        RECT 1.347 1.209 1.389 1.251 ;
        RECT 1.651 1.209 1.693 1.251 ;
        RECT 1.955 1.209 1.997 1.251 ;
        RECT 0.283 1.301 0.325 1.343 ;
        RECT 1.347 1.301 1.389 1.343 ;
        RECT 1.651 1.301 1.693 1.343 ;
        RECT 1.955 1.301 1.997 1.343 ;
        RECT 0.283 1.395 0.325 1.437 ;
        RECT 1.347 1.395 1.389 1.437 ;
        RECT 1.651 1.395 1.693 1.437 ;
        RECT 1.955 1.395 1.997 1.437 ;
        RECT 0.283 1.487 0.325 1.529 ;
        RECT 1.347 1.487 1.389 1.529 ;
        RECT 1.651 1.487 1.693 1.529 ;
        RECT 1.955 1.487 1.997 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 2.28 1.702 ;
        RECT 0.279 0.818 0.329 1.642 ;
        RECT 1.039 1.065 1.089 1.642 ;
        RECT 1.343 0.912 1.393 1.642 ;
        RECT 1.647 0.912 1.697 1.642 ;
        RECT 1.951 0.911 2.001 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 1.043 0.141 1.085 0.183 ;
        RECT 1.347 0.148 1.389 0.19 ;
        RECT 1.651 0.148 1.693 0.19 ;
        RECT 1.955 0.148 1.997 0.19 ;
        RECT 0.435 0.179 0.477 0.221 ;
        RECT 0.739 0.179 0.781 0.221 ;
        RECT 1.347 0.24 1.389 0.282 ;
        RECT 1.651 0.242 1.693 0.284 ;
        RECT 1.955 0.242 1.997 0.284 ;
        RECT 1.347 0.332 1.389 0.374 ;
        RECT 1.651 0.334 1.693 0.376 ;
        RECT 1.955 0.334 1.997 0.376 ;
      LAYER M1 ;
        RECT 1.647 0.03 1.697 0.396 ;
        RECT 1.951 0.03 2.001 0.396 ;
        RECT 1.343 0.03 1.393 0.394 ;
        RECT 0.431 0.03 0.481 0.241 ;
        RECT 0.735 0.03 0.785 0.241 ;
        RECT 1.039 0.03 1.089 0.203 ;
        RECT 0 -0.03 2.28 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 1.499 0.809 1.541 0.851 ;
      RECT 1.119 0.67 1.161 0.712 ;
      RECT 1.195 0.245 1.237 0.287 ;
      RECT 1.195 0.151 1.237 0.193 ;
      RECT 1.195 0.989 1.237 1.031 ;
      RECT 1.195 0.897 1.237 0.939 ;
      RECT 1.195 0.803 1.237 0.845 ;
      RECT 1.727 0.67 1.769 0.712 ;
      RECT 1.499 0.334 1.541 0.376 ;
      RECT 1.499 0.242 1.541 0.284 ;
      RECT 1.499 0.148 1.541 0.19 ;
      RECT 1.499 0.427 1.541 0.469 ;
      RECT 1.499 1.458 1.541 1.5 ;
      RECT 1.499 1.366 1.541 1.408 ;
      RECT 1.423 0.667 1.465 0.709 ;
      RECT 1.499 1.272 1.541 1.314 ;
      RECT 1.499 1.18 1.541 1.222 ;
      RECT 1.499 1.087 1.541 1.129 ;
      RECT 1.499 0.995 1.541 1.037 ;
      RECT 1.499 0.901 1.541 0.943 ;
      RECT 0.891 0.23 0.933 0.272 ;
      RECT 0.283 0.23 0.325 0.272 ;
      RECT 1.879 0.67 1.921 0.712 ;
      RECT 0.891 1.458 0.933 1.5 ;
      RECT 0.891 1.366 0.933 1.408 ;
      RECT 0.891 1.272 0.933 1.314 ;
      RECT 0.891 1.18 0.933 1.222 ;
      RECT 0.891 1.087 0.933 1.129 ;
      RECT 0.587 0.23 0.629 0.272 ;
      RECT 0.891 0.995 0.933 1.037 ;
    LAYER M1 ;
      RECT 1.029 0.666 1.181 0.716 ;
      RECT 1.029 0.341 1.079 0.666 ;
      RECT 0.279 0.291 1.079 0.341 ;
      RECT 1.029 0.716 1.079 0.927 ;
      RECT 0.887 0.927 1.079 0.977 ;
      RECT 0.887 0.209 0.937 0.291 ;
      RECT 0.887 0.977 0.937 1.535 ;
      RECT 0.279 0.21 0.329 0.291 ;
      RECT 0.583 0.21 0.633 0.291 ;
      RECT 1.34 0.663 1.485 0.713 ;
      RECT 1.34 0.552 1.39 0.663 ;
      RECT 1.191 0.502 1.39 0.552 ;
      RECT 1.34 0.713 1.39 0.803 ;
      RECT 1.191 0.803 1.39 0.853 ;
      RECT 1.191 0.853 1.241 1.051 ;
      RECT 1.191 0.783 1.241 0.803 ;
      RECT 1.191 0.131 1.241 0.502 ;
      RECT 1.618 0.666 1.941 0.716 ;
      RECT 1.618 0.553 1.668 0.666 ;
      RECT 1.495 0.503 1.668 0.553 ;
      RECT 1.618 0.716 1.668 0.803 ;
      RECT 1.495 0.803 1.668 0.853 ;
      RECT 1.495 0.853 1.545 1.535 ;
      RECT 1.495 0.789 1.545 0.803 ;
      RECT 1.495 0.128 1.545 0.503 ;
    LAYER PO ;
      RECT 1.733 0.071 1.763 1.612 ;
      RECT 1.885 0.071 1.915 1.612 ;
      RECT 2.037 0.071 2.067 1.612 ;
      RECT 1.581 0.071 1.611 1.612 ;
      RECT 1.125 0.071 1.155 1.612 ;
      RECT 1.277 0.071 1.307 1.612 ;
      RECT 1.429 0.071 1.459 1.61 ;
      RECT 0.973 0.072 1.003 1.61 ;
      RECT 0.061 0.072 0.091 1.61 ;
      RECT 2.189 0.072 2.219 1.61 ;
      RECT 0.821 0.072 0.851 1.61 ;
      RECT 0.213 0.072 0.243 1.61 ;
      RECT 0.669 0.072 0.699 1.61 ;
      RECT 0.365 0.072 0.395 1.61 ;
      RECT 0.517 0.072 0.547 1.61 ;
    LAYER NWELL ;
      RECT -0.115 0.679 2.395 1.801 ;
  END
END OR4X2_RVT

MACRO LATCHX1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.04 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 1.514 0.401 1.556 ;
      LAYER M1 ;
        RECT 0.355 1.423 0.405 1.576 ;
        RECT 0.249 1.313 0.405 1.423 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0342 ;
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.967 0.668 1.009 0.71 ;
      LAYER M1 ;
        RECT 0.947 0.666 1.119 0.815 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 2.715 0.158 2.757 0.2 ;
        RECT 2.715 1.3 2.757 1.342 ;
        RECT 2.715 1.392 2.757 1.434 ;
        RECT 2.715 1.484 2.757 1.526 ;
      LAYER M1 ;
        RECT 2.711 1.271 2.761 1.546 ;
        RECT 2.711 1.221 2.944 1.271 ;
        RECT 2.833 1.161 2.944 1.221 ;
        RECT 2.893 0.204 2.943 1.161 ;
        RECT 2.695 0.154 2.943 0.204 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 2.411 0.195 2.453 0.237 ;
        RECT 2.411 0.287 2.453 0.329 ;
        RECT 2.411 1.116 2.453 1.158 ;
        RECT 2.411 1.208 2.453 1.25 ;
        RECT 2.411 1.3 2.453 1.342 ;
        RECT 2.411 1.392 2.453 1.434 ;
        RECT 2.411 1.484 2.453 1.526 ;
      LAYER M1 ;
        RECT 2.407 1.119 2.457 1.546 ;
        RECT 2.407 1.069 2.791 1.119 ;
        RECT 2.681 1.009 2.791 1.069 ;
        RECT 2.741 0.359 2.791 1.009 ;
        RECT 2.407 0.309 2.791 0.359 ;
        RECT 2.407 0.148 2.457 0.309 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.435 0.881 0.477 0.923 ;
        RECT 0.587 0.895 0.629 0.937 ;
        RECT 0.435 0.973 0.477 1.015 ;
        RECT 0.587 0.987 0.629 1.029 ;
        RECT 0.435 1.065 0.477 1.107 ;
        RECT 0.587 1.079 0.629 1.121 ;
        RECT 0.891 1.097 0.933 1.139 ;
        RECT 2.259 1.122 2.301 1.164 ;
        RECT 0.891 1.189 0.933 1.231 ;
        RECT 2.563 1.208 2.605 1.25 ;
        RECT 1.499 1.212 1.541 1.254 ;
        RECT 2.259 1.214 2.301 1.256 ;
        RECT 0.891 1.281 0.933 1.323 ;
        RECT 2.563 1.3 2.605 1.342 ;
        RECT 1.499 1.304 1.541 1.346 ;
        RECT 2.259 1.306 2.301 1.348 ;
        RECT 2.563 1.392 2.605 1.434 ;
        RECT 1.499 1.396 1.541 1.438 ;
        RECT 2.259 1.398 2.301 1.44 ;
        RECT 2.563 1.484 2.605 1.526 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 3.04 1.702 ;
        RECT 1.662 1.471 1.712 1.642 ;
        RECT 1.495 1.421 1.712 1.471 ;
        RECT 2.559 1.17 2.609 1.642 ;
        RECT 1.495 1.192 1.545 1.421 ;
        RECT 0.543 1.127 0.593 1.642 ;
        RECT 2.255 1.084 2.305 1.642 ;
        RECT 0.887 1.127 0.937 1.343 ;
        RECT 0.431 1.077 0.937 1.127 ;
        RECT 0.431 0.861 0.481 1.077 ;
        RECT 0.583 0.874 0.633 1.077 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 2.563 0.158 2.605 0.2 ;
        RECT 0.435 0.2 0.477 0.242 ;
        RECT 0.587 0.2 0.629 0.242 ;
        RECT 0.435 0.292 0.477 0.334 ;
        RECT 0.587 0.292 0.629 0.334 ;
        RECT 2.259 0.292 2.301 0.334 ;
        RECT 1.499 0.308 1.541 0.35 ;
        RECT 0.891 0.324 0.933 0.366 ;
        RECT 0.435 0.388 0.477 0.43 ;
        RECT 0.587 0.388 0.629 0.43 ;
        RECT 0.891 0.416 0.933 0.458 ;
      LAYER M1 ;
        RECT 0.887 0.354 0.937 0.478 ;
        RECT 0.887 0.304 2.305 0.354 ;
        RECT 0.431 0.03 0.481 0.45 ;
        RECT 0.583 0.03 0.633 0.45 ;
        RECT 2.255 0.03 2.305 0.304 ;
        RECT 2.559 0.03 2.609 0.22 ;
        RECT 0 -0.03 3.04 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 1.879 0.2 1.921 0.242 ;
      RECT 0.283 0.852 0.325 0.894 ;
      RECT 1.423 0.2 1.465 0.242 ;
      RECT 1.347 0.914 1.389 0.956 ;
      RECT 1.803 1.14 1.845 1.182 ;
      RECT 1.347 0.43 1.389 0.472 ;
      RECT 1.803 1.048 1.845 1.09 ;
      RECT 2.107 0.53 2.149 0.572 ;
      RECT 1.043 1.291 1.085 1.333 ;
      RECT 1.043 1.199 1.085 1.241 ;
      RECT 0.283 0.245 0.325 0.287 ;
      RECT 0.739 0.414 0.781 0.456 ;
      RECT 0.739 0.506 0.781 0.548 ;
      RECT 0.663 0.622 0.705 0.664 ;
      RECT 1.195 0.438 1.237 0.48 ;
      RECT 1.347 1.006 1.389 1.048 ;
      RECT 1.195 1.042 1.237 1.084 ;
      RECT 0.739 0.76 0.781 0.802 ;
      RECT 1.651 0.912 1.693 0.954 ;
      RECT 2.487 0.664 2.529 0.706 ;
      RECT 1.195 0.53 1.237 0.572 ;
      RECT 0.283 0.521 0.325 0.563 ;
      RECT 0.283 0.429 0.325 0.471 ;
      RECT 0.283 0.337 0.325 0.379 ;
      RECT 2.107 0.812 2.149 0.854 ;
      RECT 1.195 0.95 1.237 0.992 ;
      RECT 1.651 0.524 1.693 0.566 ;
      RECT 1.955 0.529 1.997 0.571 ;
      RECT 1.955 0.812 1.997 0.854 ;
      RECT 1.271 1.53 1.313 1.572 ;
      RECT 0.283 0.944 0.325 0.986 ;
      RECT 2.183 0.664 2.225 0.706 ;
      RECT 1.271 0.1 1.313 0.142 ;
      RECT 2.031 0.1 2.073 0.142 ;
      RECT 1.575 0.622 1.617 0.664 ;
      RECT 2.639 0.608 2.681 0.65 ;
      RECT 1.879 1.53 1.921 1.572 ;
      RECT 1.803 0.414 1.845 0.456 ;
      RECT 2.031 1.53 2.073 1.572 ;
      RECT 1.195 0.858 1.237 0.9 ;
      RECT 0.283 0.76 0.325 0.802 ;
      RECT 0.283 1.036 0.325 1.078 ;
      RECT 1.347 0.522 1.389 0.564 ;
      RECT 0.739 0.852 0.781 0.894 ;
      RECT 0.739 0.322 0.781 0.364 ;
      RECT 1.043 0.422 1.085 0.464 ;
      RECT 0.663 1.53 0.705 1.572 ;
      RECT 1.423 1.53 1.465 1.572 ;
      RECT 0.739 0.226 0.781 0.268 ;
      RECT 1.347 0.822 1.389 0.864 ;
    LAYER M1 ;
      RECT 2.163 0.66 2.549 0.71 ;
      RECT 1.631 0.908 2.303 0.958 ;
      RECT 1.631 0.518 1.739 0.568 ;
      RECT 2.253 0.71 2.303 0.908 ;
      RECT 1.689 0.568 1.739 0.908 ;
      RECT 1.343 0.41 2.685 0.46 ;
      RECT 2.635 0.46 2.685 0.67 ;
      RECT 1.343 0.46 1.393 1.028 ;
      RECT 1.498 0.618 1.639 0.668 ;
      RECT 1.343 1.028 1.849 1.078 ;
      RECT 1.498 0.46 1.548 0.618 ;
      RECT 1.799 1.078 1.849 1.202 ;
      RECT 0.735 0.096 2.093 0.146 ;
      RECT 0.735 0.518 0.825 0.568 ;
      RECT 0.735 0.718 0.825 0.768 ;
      RECT 0.735 0.768 0.785 0.914 ;
      RECT 0.735 0.146 0.785 0.518 ;
      RECT 0.775 0.568 0.825 0.718 ;
      RECT 0.279 0.618 0.725 0.668 ;
      RECT 0.279 0.668 0.329 1.135 ;
      RECT 0.279 0.225 0.329 0.618 ;
      RECT 1.039 1.308 1.241 1.358 ;
      RECT 1.023 0.418 1.241 0.468 ;
      RECT 1.039 1.166 1.089 1.308 ;
      RECT 1.191 0.468 1.241 1.308 ;
      RECT 0.643 1.526 1.485 1.576 ;
      RECT 1.935 0.808 2.182 0.858 ;
      RECT 1.935 0.525 2.169 0.575 ;
      RECT 1.935 0.575 1.985 0.808 ;
      RECT 1.403 0.196 1.941 0.246 ;
      RECT 1.858 1.526 2.093 1.576 ;
    LAYER PO ;
      RECT 0.213 0.068 0.243 1.606 ;
      RECT 2.493 0.068 2.523 1.606 ;
      RECT 0.669 0.068 0.699 1.606 ;
      RECT 1.581 0.068 1.611 1.606 ;
      RECT 2.037 0.068 2.067 1.606 ;
      RECT 2.645 0.068 2.675 1.606 ;
      RECT 1.733 0.068 1.763 1.606 ;
      RECT 1.125 0.068 1.155 1.606 ;
      RECT 1.429 0.068 1.459 1.606 ;
      RECT 0.517 0.068 0.547 1.606 ;
      RECT 0.973 0.068 1.003 1.606 ;
      RECT 0.365 0.068 0.395 1.606 ;
      RECT 2.797 0.068 2.827 1.606 ;
      RECT 2.189 0.068 2.219 1.606 ;
      RECT 0.821 0.068 0.851 1.606 ;
      RECT 1.277 0.068 1.307 0.642 ;
      RECT 0.061 0.068 0.091 1.606 ;
      RECT 1.277 0.742 1.307 1.606 ;
      RECT 2.341 0.068 2.371 1.606 ;
      RECT 1.885 0.742 1.915 1.606 ;
      RECT 2.949 0.068 2.979 1.606 ;
      RECT 1.885 0.068 1.915 0.642 ;
    LAYER NWELL ;
      RECT -0.115 0.679 3.155 1.773 ;
      RECT 0.228 0.669 0.532 0.679 ;
  END
END LATCHX1_RVT

MACRO HADDX1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.75 0.401 0.792 ;
        RECT 0.967 0.75 1.009 0.792 ;
      LAYER M1 ;
        RECT 0.249 0.796 0.367 0.815 ;
        RECT 0.249 0.746 1.029 0.796 ;
        RECT 0.249 0.705 0.367 0.746 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0513 ;
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.591 0.553 0.633 ;
        RECT 1.119 0.591 1.161 0.633 ;
      LAYER M1 ;
        RECT 0.507 0.643 1.165 0.693 ;
        RECT 0.507 0.555 0.557 0.643 ;
        RECT 0.649 0.553 0.815 0.643 ;
        RECT 1.115 0.555 1.165 0.643 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0513 ;
  END B0
  PIN C1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.347 0.499 1.389 0.541 ;
        RECT 1.347 1.042 1.389 1.084 ;
      LAYER M1 ;
        RECT 1.315 1.009 1.575 1.119 ;
        RECT 1.315 0.561 1.365 1.009 ;
        RECT 1.315 0.474 1.393 0.561 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END C1
  PIN SO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.651 0.141 1.693 0.183 ;
        RECT 1.651 0.921 1.693 0.963 ;
      LAYER M1 ;
        RECT 1.631 0.917 1.879 0.967 ;
        RECT 1.671 0.857 1.879 0.917 ;
        RECT 1.671 0.187 1.721 0.857 ;
        RECT 1.631 0.137 1.721 0.187 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.343 0.325 1.385 ;
        RECT 0.739 1.343 0.781 1.385 ;
        RECT 1.043 1.343 1.085 1.385 ;
        RECT 1.499 1.39 1.541 1.432 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.976 1.702 ;
        RECT 0.279 1.323 0.329 1.642 ;
        RECT 0.735 1.323 0.785 1.642 ;
        RECT 1.039 1.318 1.089 1.642 ;
        RECT 1.495 1.363 1.545 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 1.499 0.141 1.541 0.183 ;
        RECT 0.739 0.192 0.781 0.234 ;
        RECT 0.891 0.192 0.933 0.234 ;
      LAYER M1 ;
        RECT 1.479 0.137 1.561 0.187 ;
        RECT 0.887 0.03 0.937 0.261 ;
        RECT 0.735 0.03 0.785 0.254 ;
        RECT 1.495 0.03 1.545 0.137 ;
        RECT 0 -0.03 1.976 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.452 0.387 1.502 0.613 ;
      RECT 1.419 0.613 1.502 0.663 ;
      RECT 1.175 0.337 1.502 0.387 ;
      RECT 0.638 0.889 0.861 0.939 ;
      RECT 0.811 0.939 0.861 1.126 ;
      RECT 1.419 0.663 1.469 0.736 ;
      RECT 0.811 1.126 1.265 1.176 ;
      RECT 1.215 1.176 1.265 1.317 ;
      RECT 1.191 1.317 1.265 1.411 ;
      RECT 1.215 0.387 1.265 1.126 ;
      RECT 0.263 0.174 0.655 0.224 ;
      RECT 1.013 0.237 1.621 0.287 ;
      RECT 1.571 0.287 1.621 0.734 ;
      RECT 0.092 0.36 1.063 0.41 ;
      RECT 1.013 0.287 1.063 0.36 ;
      RECT 0.092 1.057 0.649 1.107 ;
      RECT 0.092 0.41 0.142 1.057 ;
    LAYER PO ;
      RECT 0.365 0.071 0.395 1.609 ;
      RECT 0.517 0.071 0.547 1.609 ;
      RECT 0.973 0.071 1.003 1.609 ;
      RECT 1.581 0.071 1.611 1.616 ;
      RECT 1.277 0.071 1.307 1.609 ;
      RECT 0.061 0.071 0.091 1.609 ;
      RECT 1.125 0.071 1.155 1.609 ;
      RECT 0.821 0.067 0.851 1.609 ;
      RECT 1.429 0.071 1.459 1.616 ;
      RECT 0.213 0.071 0.243 1.609 ;
      RECT 0.669 0.071 0.699 1.609 ;
      RECT 1.885 0.071 1.915 1.609 ;
      RECT 1.733 0.071 1.763 1.609 ;
    LAYER CO ;
      RECT 0.587 1.061 0.629 1.103 ;
      RECT 0.283 0.179 0.325 0.221 ;
      RECT 1.423 0.655 1.465 0.697 ;
      RECT 0.663 0.893 0.705 0.935 ;
      RECT 0.891 1.13 0.933 1.172 ;
      RECT 0.587 0.178 0.629 0.22 ;
      RECT 1.195 1.343 1.237 1.385 ;
      RECT 1.575 0.617 1.617 0.659 ;
      RECT 1.195 0.341 1.237 0.383 ;
      RECT 0.435 0.364 0.477 0.406 ;
    LAYER NWELL ;
      RECT -0.115 0.679 2.091 1.773 ;
  END
END HADDX1_RVT

MACRO HEADX32_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 6.688 BY 3.344 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.119 0.679 1.161 0.721 ;
        RECT 1.271 0.679 1.313 0.721 ;
        RECT 1.423 0.679 1.465 0.721 ;
        RECT 1.575 0.679 1.617 0.721 ;
        RECT 1.727 0.679 1.769 0.721 ;
        RECT 1.879 0.679 1.921 0.721 ;
        RECT 2.031 0.679 2.073 0.721 ;
        RECT 2.183 0.679 2.225 0.721 ;
        RECT 2.335 0.679 2.377 0.721 ;
        RECT 2.487 0.679 2.529 0.721 ;
        RECT 2.639 0.679 2.681 0.721 ;
        RECT 2.791 0.679 2.833 0.721 ;
        RECT 2.943 0.679 2.985 0.721 ;
        RECT 3.095 0.679 3.137 0.721 ;
        RECT 3.247 0.679 3.289 0.721 ;
        RECT 3.399 0.679 3.441 0.721 ;
        RECT 3.551 0.679 3.593 0.721 ;
        RECT 3.703 0.679 3.745 0.721 ;
        RECT 3.855 0.679 3.897 0.721 ;
        RECT 4.007 0.679 4.049 0.721 ;
        RECT 4.159 0.679 4.201 0.721 ;
        RECT 4.311 0.679 4.353 0.721 ;
        RECT 4.463 0.679 4.505 0.721 ;
        RECT 4.615 0.679 4.657 0.721 ;
        RECT 4.767 0.679 4.809 0.721 ;
        RECT 4.919 0.679 4.961 0.721 ;
        RECT 5.071 0.679 5.113 0.721 ;
        RECT 5.223 0.679 5.265 0.721 ;
        RECT 5.375 0.679 5.417 0.721 ;
        RECT 5.527 0.679 5.569 0.721 ;
        RECT 5.679 0.679 5.721 0.721 ;
        RECT 5.831 0.679 5.873 0.721 ;
      LAYER M1 ;
        RECT 1.099 0.67 5.893 0.73 ;
        RECT 1.12 0.553 1.31 0.67 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0 ;
  END SLEEP
  PIN VDD
    DIRECTION OUTPUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 5.907 0.853 5.949 0.895 ;
        RECT 5.907 0.945 5.949 0.987 ;
        RECT 1.043 1.037 1.085 1.079 ;
        RECT 1.347 1.037 1.389 1.079 ;
        RECT 1.651 1.037 1.693 1.079 ;
        RECT 1.955 1.037 1.997 1.079 ;
        RECT 2.259 1.037 2.301 1.079 ;
        RECT 2.563 1.037 2.605 1.079 ;
        RECT 2.867 1.037 2.909 1.079 ;
        RECT 3.171 1.037 3.213 1.079 ;
        RECT 3.475 1.037 3.517 1.079 ;
        RECT 3.779 1.037 3.821 1.079 ;
        RECT 4.083 1.037 4.125 1.079 ;
        RECT 4.387 1.037 4.429 1.079 ;
        RECT 4.691 1.037 4.733 1.079 ;
        RECT 4.995 1.037 5.037 1.079 ;
        RECT 5.299 1.037 5.341 1.079 ;
        RECT 5.603 1.037 5.645 1.079 ;
        RECT 5.907 1.037 5.949 1.079 ;
        RECT 1.043 1.129 1.085 1.171 ;
        RECT 1.347 1.129 1.389 1.171 ;
        RECT 1.651 1.129 1.693 1.171 ;
        RECT 1.955 1.129 1.997 1.171 ;
        RECT 2.259 1.129 2.301 1.171 ;
        RECT 2.563 1.129 2.605 1.171 ;
        RECT 2.867 1.129 2.909 1.171 ;
        RECT 3.171 1.129 3.213 1.171 ;
        RECT 3.475 1.129 3.517 1.171 ;
        RECT 3.779 1.129 3.821 1.171 ;
        RECT 4.083 1.129 4.125 1.171 ;
        RECT 4.387 1.129 4.429 1.171 ;
        RECT 4.691 1.129 4.733 1.171 ;
        RECT 4.995 1.129 5.037 1.171 ;
        RECT 5.299 1.129 5.341 1.171 ;
        RECT 5.603 1.129 5.645 1.171 ;
        RECT 5.907 1.129 5.949 1.171 ;
        RECT 1.043 1.221 1.085 1.263 ;
        RECT 1.347 1.221 1.389 1.263 ;
        RECT 1.651 1.221 1.693 1.263 ;
        RECT 1.955 1.221 1.997 1.263 ;
        RECT 2.259 1.221 2.301 1.263 ;
        RECT 2.563 1.221 2.605 1.263 ;
        RECT 2.867 1.221 2.909 1.263 ;
        RECT 3.171 1.221 3.213 1.263 ;
        RECT 3.475 1.221 3.517 1.263 ;
        RECT 3.779 1.221 3.821 1.263 ;
        RECT 4.083 1.221 4.125 1.263 ;
        RECT 4.387 1.221 4.429 1.263 ;
        RECT 4.691 1.221 4.733 1.263 ;
        RECT 4.995 1.221 5.037 1.263 ;
        RECT 5.299 1.221 5.341 1.263 ;
        RECT 5.603 1.221 5.645 1.263 ;
        RECT 5.907 1.221 5.949 1.263 ;
        RECT 1.043 1.313 1.085 1.355 ;
        RECT 1.347 1.313 1.389 1.355 ;
        RECT 1.651 1.313 1.693 1.355 ;
        RECT 1.955 1.313 1.997 1.355 ;
        RECT 2.259 1.313 2.301 1.355 ;
        RECT 2.563 1.313 2.605 1.355 ;
        RECT 2.867 1.313 2.909 1.355 ;
        RECT 3.171 1.313 3.213 1.355 ;
        RECT 3.475 1.313 3.517 1.355 ;
        RECT 3.779 1.313 3.821 1.355 ;
        RECT 4.083 1.313 4.125 1.355 ;
        RECT 4.387 1.313 4.429 1.355 ;
        RECT 4.691 1.313 4.733 1.355 ;
        RECT 4.995 1.313 5.037 1.355 ;
        RECT 5.299 1.313 5.341 1.355 ;
        RECT 5.603 1.313 5.645 1.355 ;
        RECT 5.907 1.313 5.949 1.355 ;
        RECT 1.043 1.407 1.085 1.449 ;
        RECT 1.347 1.407 1.389 1.449 ;
        RECT 1.651 1.407 1.693 1.449 ;
        RECT 1.955 1.407 1.997 1.449 ;
        RECT 2.259 1.407 2.301 1.449 ;
        RECT 2.563 1.407 2.605 1.449 ;
        RECT 2.867 1.407 2.909 1.449 ;
        RECT 3.171 1.407 3.213 1.449 ;
        RECT 3.475 1.407 3.517 1.449 ;
        RECT 3.779 1.407 3.821 1.449 ;
        RECT 4.083 1.407 4.125 1.449 ;
        RECT 4.387 1.407 4.429 1.449 ;
        RECT 4.691 1.407 4.733 1.449 ;
        RECT 4.995 1.407 5.037 1.449 ;
        RECT 5.299 1.407 5.341 1.449 ;
        RECT 5.603 1.407 5.645 1.449 ;
        RECT 5.907 1.407 5.949 1.449 ;
        RECT 1.043 1.499 1.085 1.541 ;
        RECT 1.347 1.499 1.389 1.541 ;
        RECT 1.651 1.499 1.693 1.541 ;
        RECT 1.955 1.499 1.997 1.541 ;
        RECT 2.259 1.499 2.301 1.541 ;
        RECT 2.563 1.499 2.605 1.541 ;
        RECT 2.867 1.499 2.909 1.541 ;
        RECT 3.171 1.499 3.213 1.541 ;
        RECT 3.475 1.499 3.517 1.541 ;
        RECT 3.779 1.499 3.821 1.541 ;
        RECT 4.083 1.499 4.125 1.541 ;
        RECT 4.387 1.499 4.429 1.541 ;
        RECT 4.691 1.499 4.733 1.541 ;
        RECT 4.995 1.499 5.037 1.541 ;
        RECT 5.299 1.499 5.341 1.541 ;
        RECT 5.603 1.499 5.645 1.541 ;
        RECT 5.907 1.499 5.949 1.541 ;
      LAYER M1 ;
        RECT 0 1.642 6.688 1.702 ;
        RECT 3.471 1.017 3.521 1.642 ;
        RECT 3.775 1.017 3.825 1.642 ;
        RECT 4.079 1.017 4.129 1.642 ;
        RECT 4.383 1.017 4.433 1.642 ;
        RECT 4.687 1.017 4.737 1.642 ;
        RECT 4.991 1.017 5.041 1.642 ;
        RECT 5.295 1.017 5.345 1.642 ;
        RECT 5.599 1.017 5.649 1.642 ;
        RECT 5.903 0.833 5.953 1.642 ;
        RECT 1.039 1.017 1.089 1.642 ;
        RECT 1.343 1.017 1.393 1.642 ;
        RECT 1.647 1.017 1.697 1.642 ;
        RECT 1.951 1.017 2.001 1.642 ;
        RECT 2.255 1.017 2.305 1.642 ;
        RECT 2.559 1.017 2.609 1.642 ;
        RECT 2.863 1.017 2.913 1.642 ;
        RECT 3.167 1.017 3.217 1.642 ;
    END
  END VDD
  PIN VDDG
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.195 0.853 1.237 0.895 ;
        RECT 1.499 0.853 1.541 0.895 ;
        RECT 1.803 0.853 1.845 0.895 ;
        RECT 2.107 0.853 2.149 0.895 ;
        RECT 2.411 0.853 2.453 0.895 ;
        RECT 2.715 0.853 2.757 0.895 ;
        RECT 3.019 0.853 3.061 0.895 ;
        RECT 3.323 0.853 3.365 0.895 ;
        RECT 3.627 0.853 3.669 0.895 ;
        RECT 3.931 0.853 3.973 0.895 ;
        RECT 4.235 0.853 4.277 0.895 ;
        RECT 4.539 0.853 4.581 0.895 ;
        RECT 4.843 0.853 4.885 0.895 ;
        RECT 5.147 0.853 5.189 0.895 ;
        RECT 5.451 0.853 5.493 0.895 ;
        RECT 5.755 0.853 5.797 0.895 ;
        RECT 1.195 0.945 1.237 0.987 ;
        RECT 1.499 0.945 1.541 0.987 ;
        RECT 1.803 0.945 1.845 0.987 ;
        RECT 2.107 0.945 2.149 0.987 ;
        RECT 2.411 0.945 2.453 0.987 ;
        RECT 2.715 0.945 2.757 0.987 ;
        RECT 3.019 0.945 3.061 0.987 ;
        RECT 3.323 0.945 3.365 0.987 ;
        RECT 3.627 0.945 3.669 0.987 ;
        RECT 3.931 0.945 3.973 0.987 ;
        RECT 4.235 0.945 4.277 0.987 ;
        RECT 4.539 0.945 4.581 0.987 ;
        RECT 4.843 0.945 4.885 0.987 ;
        RECT 5.147 0.945 5.189 0.987 ;
        RECT 5.451 0.945 5.493 0.987 ;
        RECT 5.755 0.945 5.797 0.987 ;
        RECT 0.739 1.011 0.781 1.053 ;
        RECT 1.195 1.037 1.237 1.079 ;
        RECT 1.499 1.037 1.541 1.079 ;
        RECT 1.803 1.037 1.845 1.079 ;
        RECT 2.107 1.037 2.149 1.079 ;
        RECT 2.411 1.037 2.453 1.079 ;
        RECT 2.715 1.037 2.757 1.079 ;
        RECT 3.019 1.037 3.061 1.079 ;
        RECT 3.323 1.037 3.365 1.079 ;
        RECT 3.627 1.037 3.669 1.079 ;
        RECT 3.931 1.037 3.973 1.079 ;
        RECT 4.235 1.037 4.277 1.079 ;
        RECT 4.539 1.037 4.581 1.079 ;
        RECT 4.843 1.037 4.885 1.079 ;
        RECT 5.147 1.037 5.189 1.079 ;
        RECT 5.451 1.037 5.493 1.079 ;
        RECT 5.755 1.037 5.797 1.079 ;
        RECT 0.739 1.103 0.781 1.145 ;
        RECT 1.195 1.129 1.237 1.171 ;
        RECT 1.499 1.129 1.541 1.171 ;
        RECT 1.803 1.129 1.845 1.171 ;
        RECT 2.107 1.129 2.149 1.171 ;
        RECT 2.411 1.129 2.453 1.171 ;
        RECT 2.715 1.129 2.757 1.171 ;
        RECT 3.019 1.129 3.061 1.171 ;
        RECT 3.323 1.129 3.365 1.171 ;
        RECT 3.627 1.129 3.669 1.171 ;
        RECT 3.931 1.129 3.973 1.171 ;
        RECT 4.235 1.129 4.277 1.171 ;
        RECT 4.539 1.129 4.581 1.171 ;
        RECT 4.843 1.129 4.885 1.171 ;
        RECT 5.147 1.129 5.189 1.171 ;
        RECT 5.451 1.129 5.493 1.171 ;
        RECT 5.755 1.129 5.797 1.171 ;
        RECT 1.195 1.221 1.237 1.263 ;
        RECT 1.499 1.221 1.541 1.263 ;
        RECT 1.803 1.221 1.845 1.263 ;
        RECT 2.107 1.221 2.149 1.263 ;
        RECT 2.411 1.221 2.453 1.263 ;
        RECT 2.715 1.221 2.757 1.263 ;
        RECT 3.019 1.221 3.061 1.263 ;
        RECT 3.323 1.221 3.365 1.263 ;
        RECT 3.627 1.221 3.669 1.263 ;
        RECT 3.931 1.221 3.973 1.263 ;
        RECT 4.235 1.221 4.277 1.263 ;
        RECT 4.539 1.221 4.581 1.263 ;
        RECT 4.843 1.221 4.885 1.263 ;
        RECT 5.147 1.221 5.189 1.263 ;
        RECT 5.451 1.221 5.493 1.263 ;
        RECT 5.755 1.221 5.797 1.263 ;
        RECT 1.195 1.313 1.237 1.355 ;
        RECT 1.499 1.313 1.541 1.355 ;
        RECT 1.803 1.313 1.845 1.355 ;
        RECT 2.107 1.313 2.149 1.355 ;
        RECT 2.411 1.313 2.453 1.355 ;
        RECT 2.715 1.313 2.757 1.355 ;
        RECT 3.019 1.313 3.061 1.355 ;
        RECT 3.323 1.313 3.365 1.355 ;
        RECT 3.627 1.313 3.669 1.355 ;
        RECT 3.931 1.313 3.973 1.355 ;
        RECT 4.235 1.313 4.277 1.355 ;
        RECT 4.539 1.313 4.581 1.355 ;
        RECT 4.843 1.313 4.885 1.355 ;
        RECT 5.147 1.313 5.189 1.355 ;
        RECT 5.451 1.313 5.493 1.355 ;
        RECT 5.755 1.313 5.797 1.355 ;
        RECT 1.195 1.407 1.237 1.449 ;
        RECT 1.499 1.407 1.541 1.449 ;
        RECT 1.803 1.407 1.845 1.449 ;
        RECT 2.107 1.407 2.149 1.449 ;
        RECT 2.411 1.407 2.453 1.449 ;
        RECT 2.715 1.407 2.757 1.449 ;
        RECT 3.019 1.407 3.061 1.449 ;
        RECT 3.323 1.407 3.365 1.449 ;
        RECT 3.627 1.407 3.669 1.449 ;
        RECT 3.931 1.407 3.973 1.449 ;
        RECT 4.235 1.407 4.277 1.449 ;
        RECT 4.539 1.407 4.581 1.449 ;
        RECT 4.843 1.407 4.885 1.449 ;
        RECT 5.147 1.407 5.189 1.449 ;
        RECT 5.451 1.407 5.493 1.449 ;
        RECT 5.755 1.407 5.797 1.449 ;
        RECT 1.195 1.499 1.237 1.541 ;
        RECT 1.499 1.499 1.541 1.541 ;
        RECT 1.803 1.499 1.845 1.541 ;
        RECT 2.107 1.499 2.149 1.541 ;
        RECT 2.411 1.499 2.453 1.541 ;
        RECT 2.715 1.499 2.757 1.541 ;
        RECT 3.019 1.499 3.061 1.541 ;
        RECT 3.323 1.499 3.365 1.541 ;
        RECT 3.627 1.499 3.669 1.541 ;
        RECT 3.931 1.499 3.973 1.541 ;
        RECT 4.235 1.499 4.277 1.541 ;
        RECT 4.539 1.499 4.581 1.541 ;
        RECT 4.843 1.499 4.885 1.541 ;
        RECT 5.147 1.499 5.189 1.541 ;
        RECT 5.451 1.499 5.493 1.541 ;
        RECT 5.755 1.499 5.797 1.541 ;
      LAYER M1 ;
        RECT 0.73 1.119 0.79 1.165 ;
        RECT 0.666 1.009 0.856 1.119 ;
        RECT 0.73 0.856 5.801 0.881 ;
        RECT 0.735 0.831 5.801 0.856 ;
        RECT 3.319 0.881 3.369 1.561 ;
        RECT 3.623 0.881 3.673 1.561 ;
        RECT 3.927 0.881 3.977 1.561 ;
        RECT 4.231 0.881 4.281 1.561 ;
        RECT 4.535 0.881 4.585 1.561 ;
        RECT 4.839 0.881 4.889 1.561 ;
        RECT 5.143 0.881 5.193 1.561 ;
        RECT 5.447 0.881 5.497 1.561 ;
        RECT 5.751 0.881 5.801 1.561 ;
        RECT 1.191 0.881 1.241 1.561 ;
        RECT 1.495 0.881 1.545 1.561 ;
        RECT 1.799 0.881 1.849 1.561 ;
        RECT 2.103 0.881 2.153 1.561 ;
        RECT 2.407 0.881 2.457 1.561 ;
        RECT 2.711 0.881 2.761 1.561 ;
        RECT 3.015 0.881 3.065 1.561 ;
        RECT 0.73 0.881 0.79 1.009 ;
    END
  END VDDG
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 3.399 -0.021 3.441 0.021 ;
        RECT 3.551 -0.021 3.593 0.021 ;
        RECT 3.703 -0.021 3.745 0.021 ;
        RECT 3.855 -0.021 3.897 0.021 ;
        RECT 4.007 -0.021 4.049 0.021 ;
        RECT 4.159 -0.021 4.201 0.021 ;
        RECT 4.311 -0.021 4.353 0.021 ;
        RECT 4.463 -0.021 4.505 0.021 ;
        RECT 4.615 -0.021 4.657 0.021 ;
        RECT 4.767 -0.021 4.809 0.021 ;
        RECT 4.919 -0.021 4.961 0.021 ;
        RECT 5.071 -0.021 5.113 0.021 ;
        RECT 5.223 -0.021 5.265 0.021 ;
        RECT 5.375 -0.021 5.417 0.021 ;
        RECT 5.527 -0.021 5.569 0.021 ;
        RECT 5.679 -0.021 5.721 0.021 ;
        RECT 5.831 -0.021 5.873 0.021 ;
        RECT 5.983 -0.021 6.025 0.021 ;
        RECT 6.135 -0.021 6.177 0.021 ;
        RECT 6.287 -0.021 6.329 0.021 ;
        RECT 6.439 -0.021 6.481 0.021 ;
        RECT 6.591 -0.021 6.633 0.021 ;
        RECT 0.055 3.323 0.097 3.365 ;
        RECT 0.207 3.323 0.249 3.365 ;
        RECT 0.359 3.323 0.401 3.365 ;
        RECT 0.511 3.323 0.553 3.365 ;
        RECT 0.663 3.323 0.705 3.365 ;
        RECT 0.815 3.323 0.857 3.365 ;
        RECT 0.967 3.323 1.009 3.365 ;
        RECT 1.119 3.323 1.161 3.365 ;
        RECT 1.271 3.323 1.313 3.365 ;
        RECT 1.423 3.323 1.465 3.365 ;
        RECT 1.575 3.323 1.617 3.365 ;
        RECT 1.727 3.323 1.769 3.365 ;
        RECT 1.879 3.323 1.921 3.365 ;
        RECT 2.031 3.323 2.073 3.365 ;
        RECT 2.183 3.323 2.225 3.365 ;
        RECT 2.335 3.323 2.377 3.365 ;
        RECT 2.487 3.323 2.529 3.365 ;
        RECT 2.639 3.323 2.681 3.365 ;
        RECT 2.791 3.323 2.833 3.365 ;
        RECT 2.943 3.323 2.985 3.365 ;
        RECT 3.095 3.323 3.137 3.365 ;
        RECT 3.247 3.323 3.289 3.365 ;
        RECT 3.399 3.323 3.441 3.365 ;
        RECT 3.551 3.323 3.593 3.365 ;
        RECT 3.703 3.323 3.745 3.365 ;
        RECT 3.855 3.323 3.897 3.365 ;
        RECT 4.007 3.323 4.049 3.365 ;
        RECT 4.159 3.323 4.201 3.365 ;
        RECT 4.311 3.323 4.353 3.365 ;
        RECT 4.463 3.323 4.505 3.365 ;
        RECT 4.615 3.323 4.657 3.365 ;
        RECT 4.767 3.323 4.809 3.365 ;
        RECT 4.919 3.323 4.961 3.365 ;
        RECT 5.071 3.323 5.113 3.365 ;
        RECT 5.223 3.323 5.265 3.365 ;
        RECT 5.375 3.323 5.417 3.365 ;
        RECT 5.527 3.323 5.569 3.365 ;
        RECT 5.679 3.323 5.721 3.365 ;
        RECT 5.831 3.323 5.873 3.365 ;
        RECT 5.983 3.323 6.025 3.365 ;
        RECT 6.135 3.323 6.177 3.365 ;
        RECT 6.287 3.323 6.329 3.365 ;
        RECT 6.439 3.323 6.481 3.365 ;
        RECT 6.591 3.323 6.633 3.365 ;
      LAYER M1 ;
        RECT 0 -0.03 6.688 0.03 ;
        RECT 0 3.314 6.688 3.374 ;
    END
  END VSS
  OBS
    LAYER PO ;
      RECT 4.165 1.739 4.195 3.252 ;
      RECT 4.317 1.739 4.347 3.252 ;
      RECT 4.469 1.739 4.499 3.252 ;
      RECT 4.621 1.739 4.651 3.252 ;
      RECT 4.773 1.739 4.803 3.252 ;
      RECT 4.925 1.739 4.955 3.252 ;
      RECT 5.077 1.739 5.107 3.252 ;
      RECT 5.229 1.739 5.259 3.252 ;
      RECT 5.381 1.739 5.411 3.252 ;
      RECT 5.533 1.739 5.563 3.252 ;
      RECT 5.685 1.739 5.715 3.252 ;
      RECT 5.989 1.739 6.019 3.252 ;
      RECT 2.037 1.739 2.067 3.252 ;
      RECT 1.885 1.739 1.915 3.252 ;
      RECT 0.669 1.739 0.699 3.252 ;
      RECT 6.597 0.108 6.627 1.621 ;
      RECT 6.445 0.108 6.475 1.621 ;
      RECT 6.293 0.108 6.323 1.621 ;
      RECT 6.141 0.108 6.171 1.621 ;
      RECT 0.517 0.107 0.547 1.62 ;
      RECT 0.365 0.107 0.395 1.62 ;
      RECT 0.213 0.107 0.243 1.62 ;
      RECT 0.061 0.107 0.091 1.62 ;
      RECT 0.517 1.739 0.547 3.252 ;
      RECT 0.365 1.739 0.395 3.252 ;
      RECT 0.213 1.739 0.243 3.252 ;
      RECT 0.061 1.739 0.091 3.252 ;
      RECT 6.597 1.739 6.627 3.252 ;
      RECT 6.445 1.739 6.475 3.252 ;
      RECT 6.293 1.739 6.323 3.252 ;
      RECT 6.141 1.739 6.171 3.252 ;
      RECT 2.645 1.739 2.675 3.252 ;
      RECT 2.493 1.739 2.523 3.252 ;
      RECT 3.557 1.739 3.587 3.252 ;
      RECT 2.341 1.739 2.371 3.252 ;
      RECT 2.189 1.739 2.219 3.252 ;
      RECT 2.797 1.739 2.827 3.252 ;
      RECT 2.949 1.739 2.979 3.252 ;
      RECT 3.101 1.739 3.131 3.252 ;
      RECT 3.253 1.739 3.283 3.252 ;
      RECT 3.405 1.739 3.435 3.252 ;
      RECT 2.645 0.108 2.675 1.621 ;
      RECT 2.493 0.108 2.523 1.621 ;
      RECT 3.557 0.108 3.587 1.621 ;
      RECT 2.341 0.108 2.371 1.621 ;
      RECT 2.189 0.108 2.219 1.621 ;
      RECT 2.037 0.108 2.067 1.621 ;
      RECT 1.885 0.108 1.915 1.621 ;
      RECT 0.669 0.108 0.699 1.621 ;
      RECT 1.581 0.108 1.611 1.621 ;
      RECT 0.821 0.108 0.851 1.621 ;
      RECT 0.973 0.108 1.003 1.621 ;
      RECT 1.429 0.108 1.459 1.621 ;
      RECT 1.733 0.108 1.763 1.621 ;
      RECT 1.125 0.108 1.155 1.621 ;
      RECT 1.277 0.108 1.307 1.621 ;
      RECT 3.709 0.108 3.739 1.621 ;
      RECT 3.861 0.108 3.891 1.621 ;
      RECT 4.013 0.108 4.043 1.621 ;
      RECT 4.165 0.108 4.195 1.621 ;
      RECT 4.317 0.108 4.347 1.621 ;
      RECT 4.469 0.108 4.499 1.621 ;
      RECT 4.621 0.108 4.651 1.621 ;
      RECT 4.773 0.108 4.803 1.621 ;
      RECT 4.925 0.108 4.955 1.621 ;
      RECT 5.077 0.108 5.107 1.621 ;
      RECT 5.229 0.108 5.259 1.621 ;
      RECT 5.381 0.108 5.411 1.621 ;
      RECT 5.533 0.108 5.563 1.621 ;
      RECT 5.685 0.108 5.715 1.621 ;
      RECT 5.837 0.108 5.867 1.621 ;
      RECT 5.989 0.108 6.019 1.621 ;
      RECT 3.405 0.108 3.435 1.621 ;
      RECT 3.253 0.108 3.283 1.621 ;
      RECT 3.101 0.108 3.131 1.621 ;
      RECT 2.949 0.108 2.979 1.621 ;
      RECT 2.797 0.108 2.827 1.621 ;
      RECT 5.837 1.739 5.867 3.252 ;
      RECT 1.581 1.739 1.611 3.252 ;
      RECT 0.821 1.739 0.851 3.252 ;
      RECT 0.973 1.739 1.003 3.252 ;
      RECT 1.429 1.739 1.459 3.252 ;
      RECT 1.733 1.739 1.763 3.252 ;
      RECT 1.125 1.739 1.155 3.252 ;
      RECT 1.277 1.739 1.307 3.252 ;
      RECT 3.709 1.739 3.739 3.252 ;
      RECT 3.861 1.739 3.891 3.252 ;
      RECT 4.013 1.739 4.043 3.252 ;
    LAYER NWELL ;
      RECT 0.571 0.679 6.109 2.665 ;
  END
END HEADX32_RVT

MACRO DELLN1X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.04 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.679 0.401 0.721 ;
      LAYER M1 ;
        RECT 0.097 0.725 0.21 0.815 ;
        RECT 0.097 0.675 0.421 0.725 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0105 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 2.411 0.151 2.453 0.193 ;
        RECT 2.715 0.151 2.757 0.193 ;
        RECT 2.411 0.243 2.453 0.285 ;
        RECT 2.715 0.243 2.757 0.285 ;
        RECT 2.411 0.335 2.453 0.377 ;
        RECT 2.715 0.335 2.757 0.377 ;
        RECT 2.411 0.427 2.453 0.469 ;
        RECT 2.715 0.427 2.757 0.469 ;
        RECT 2.411 1.027 2.453 1.069 ;
        RECT 2.715 1.027 2.757 1.069 ;
        RECT 2.411 1.119 2.453 1.161 ;
        RECT 2.715 1.119 2.757 1.161 ;
        RECT 2.411 1.211 2.453 1.253 ;
        RECT 2.715 1.211 2.757 1.253 ;
        RECT 2.411 1.303 2.453 1.345 ;
        RECT 2.715 1.303 2.757 1.345 ;
        RECT 2.411 1.395 2.453 1.437 ;
        RECT 2.715 1.395 2.757 1.437 ;
        RECT 2.411 1.487 2.453 1.529 ;
        RECT 2.715 1.487 2.757 1.529 ;
      LAYER M1 ;
        RECT 2.407 0.942 2.457 1.549 ;
        RECT 2.711 0.942 2.761 1.549 ;
        RECT 2.407 0.892 2.801 0.942 ;
        RECT 2.751 0.663 2.801 0.892 ;
        RECT 2.751 0.587 2.943 0.663 ;
        RECT 2.407 0.537 2.943 0.587 ;
        RECT 2.407 0.131 2.457 0.537 ;
        RECT 2.711 0.131 2.761 0.537 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.663 0.573 0.705 0.615 ;
        RECT 0.815 0.573 0.857 0.615 ;
        RECT 1.575 0.603 1.617 0.645 ;
        RECT 1.727 0.603 1.769 0.645 ;
        RECT 1.195 0.817 1.237 0.859 ;
        RECT 2.107 0.836 2.149 0.878 ;
        RECT 0.283 0.837 0.325 0.879 ;
        RECT 1.195 0.909 1.237 0.951 ;
        RECT 2.107 0.928 2.149 0.97 ;
        RECT 0.283 0.929 0.325 0.971 ;
        RECT 2.107 1.02 2.149 1.062 ;
        RECT 2.563 1.027 2.605 1.069 ;
        RECT 2.107 1.112 2.149 1.154 ;
        RECT 2.563 1.119 2.605 1.161 ;
        RECT 2.107 1.204 2.149 1.246 ;
        RECT 1.499 1.208 1.541 1.25 ;
        RECT 2.563 1.211 2.605 1.253 ;
        RECT 0.587 1.292 0.629 1.334 ;
        RECT 1.499 1.3 1.541 1.342 ;
        RECT 2.563 1.303 2.605 1.345 ;
        RECT 0.587 1.384 0.629 1.426 ;
        RECT 1.499 1.392 1.541 1.434 ;
        RECT 2.563 1.395 2.605 1.437 ;
        RECT 0.587 1.476 0.629 1.518 ;
        RECT 1.499 1.484 1.541 1.526 ;
        RECT 2.563 1.487 2.605 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 3.04 1.702 ;
        RECT 0.583 1.29 0.633 1.642 ;
        RECT 0.543 1.24 0.633 1.29 ;
        RECT 1.495 1.15 1.545 1.642 ;
        RECT 1.455 1.1 1.545 1.15 ;
        RECT 0.543 1.09 0.593 1.24 ;
        RECT 2.559 0.992 2.609 1.642 ;
        RECT 0.543 1.04 0.621 1.09 ;
        RECT 1.455 0.95 1.505 1.1 ;
        RECT 0.279 0.817 0.329 1.642 ;
        RECT 1.191 0.797 1.241 1.642 ;
        RECT 2.103 0.816 2.153 1.642 ;
        RECT 1.455 0.9 1.549 0.95 ;
        RECT 1.499 0.649 1.549 0.9 ;
        RECT 0.571 0.619 0.621 1.04 ;
        RECT 1.499 0.599 1.789 0.649 ;
        RECT 0.571 0.569 0.877 0.619 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 2.563 0.149 2.605 0.191 ;
        RECT 2.563 0.241 2.605 0.283 ;
        RECT 2.107 0.301 2.149 0.343 ;
        RECT 2.563 0.333 2.605 0.375 ;
        RECT 0.587 0.371 0.629 0.413 ;
        RECT 1.499 0.381 1.541 0.423 ;
        RECT 2.107 0.393 2.149 0.435 ;
        RECT 1.499 0.474 1.541 0.516 ;
        RECT 0.283 0.478 0.325 0.52 ;
        RECT 2.107 0.485 2.149 0.527 ;
        RECT 1.195 0.488 1.237 0.53 ;
        RECT 1.575 1.004 1.617 1.046 ;
        RECT 1.727 1.004 1.769 1.046 ;
        RECT 0.663 1.144 0.705 1.186 ;
        RECT 0.815 1.144 0.857 1.186 ;
      LAYER M1 ;
        RECT 0.643 1.14 0.977 1.19 ;
        RECT 1.555 1 1.889 1.05 ;
        RECT 1.839 0.549 1.889 1 ;
        RECT 0.927 0.519 0.977 1.14 ;
        RECT 1.495 0.499 1.889 0.549 ;
        RECT 0.583 0.469 0.977 0.519 ;
        RECT 1.495 0.248 1.545 0.499 ;
        RECT 0.583 0.248 0.633 0.469 ;
        RECT 0.583 0.198 1.129 0.248 ;
        RECT 1.495 0.198 2.041 0.248 ;
        RECT 1.191 0.03 1.241 0.55 ;
        RECT 2.103 0.03 2.153 0.547 ;
        RECT 0.279 0.03 0.329 0.54 ;
        RECT 2.559 0.03 2.609 0.41 ;
        RECT 1.079 0.03 1.129 0.198 ;
        RECT 1.991 0.03 2.041 0.198 ;
        RECT 0 -0.03 3.04 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 1.955 1.291 1.997 1.333 ;
      RECT 1.879 0.1 1.921 0.142 ;
      RECT 1.955 1.475 1.997 1.517 ;
      RECT 1.955 1.198 1.997 1.24 ;
      RECT 1.043 0.367 1.085 0.409 ;
      RECT 1.955 1.106 1.997 1.148 ;
      RECT 1.955 1.106 1.997 1.148 ;
      RECT 1.955 1.198 1.997 1.24 ;
      RECT 2.259 1.206 2.301 1.248 ;
      RECT 1.955 0.391 1.997 0.433 ;
      RECT 1.955 0.391 1.997 0.433 ;
      RECT 2.259 0.301 2.301 0.343 ;
      RECT 2.183 0.664 2.225 0.706 ;
      RECT 2.259 0.93 2.301 0.972 ;
      RECT 2.259 1.206 2.301 1.248 ;
      RECT 2.487 0.664 2.529 0.706 ;
      RECT 2.259 1.114 2.301 1.156 ;
      RECT 1.347 0.817 1.389 0.859 ;
      RECT 1.347 0.817 1.389 0.859 ;
      RECT 1.347 0.909 1.389 0.951 ;
      RECT 1.347 0.909 1.389 0.951 ;
      RECT 0.435 0.837 0.477 0.879 ;
      RECT 0.435 0.837 0.477 0.879 ;
      RECT 0.435 0.929 0.477 0.971 ;
      RECT 1.955 1.291 1.997 1.333 ;
      RECT 0.435 0.929 0.477 0.971 ;
      RECT 1.043 1.379 1.085 1.421 ;
      RECT 0.435 0.498 0.477 0.54 ;
      RECT 1.043 0.367 1.085 0.409 ;
      RECT 1.043 1.287 1.085 1.329 ;
      RECT 1.043 1.287 1.085 1.329 ;
      RECT 1.043 1.379 1.085 1.421 ;
      RECT 0.435 0.498 0.477 0.54 ;
      RECT 1.955 1.383 1.997 1.425 ;
      RECT 0.967 0.1 1.009 0.142 ;
      RECT 2.259 1.022 2.301 1.064 ;
      RECT 2.259 0.93 2.301 0.972 ;
      RECT 2.259 0.485 2.301 0.527 ;
      RECT 2.259 0.393 2.301 0.435 ;
      RECT 2.259 0.393 2.301 0.435 ;
      RECT 2.639 0.664 2.681 0.706 ;
      RECT 2.259 1.022 2.301 1.064 ;
      RECT 2.259 1.114 2.301 1.156 ;
      RECT 1.955 1.383 1.997 1.425 ;
      RECT 1.955 0.483 1.997 0.525 ;
      RECT 1.043 0.459 1.085 0.501 ;
      RECT 1.955 1.475 1.997 1.517 ;
      RECT 1.043 1.472 1.085 1.514 ;
      RECT 1.043 1.472 1.085 1.514 ;
      RECT 1.347 0.488 1.389 0.53 ;
      RECT 1.271 0.679 1.313 0.721 ;
      RECT 1.043 0.459 1.085 0.501 ;
    LAYER M1 ;
      RECT 1.039 0.675 1.333 0.725 ;
      RECT 1.039 0.725 1.089 1.534 ;
      RECT 1.039 0.347 1.089 0.675 ;
      RECT 0.431 0.096 1.029 0.146 ;
      RECT 0.431 0.541 0.521 0.591 ;
      RECT 0.431 0.825 0.481 0.999 ;
      RECT 0.431 0.146 0.481 0.541 ;
      RECT 0.431 0.775 0.521 0.825 ;
      RECT 0.471 0.591 0.521 0.775 ;
      RECT 1.951 0.66 2.245 0.71 ;
      RECT 1.951 0.71 2.001 1.537 ;
      RECT 1.951 0.371 2.001 0.66 ;
      RECT 1.343 0.096 1.941 0.146 ;
      RECT 1.343 0.146 1.393 0.532 ;
      RECT 1.343 0.775 1.433 0.825 ;
      RECT 1.343 0.825 1.393 0.971 ;
      RECT 1.383 0.582 1.433 0.775 ;
      RECT 1.343 0.532 1.433 0.582 ;
      RECT 2.295 0.66 2.701 0.71 ;
      RECT 2.255 0.937 2.305 1.269 ;
      RECT 2.255 0.887 2.345 0.937 ;
      RECT 2.295 0.71 2.345 0.887 ;
      RECT 2.255 0.281 2.305 0.532 ;
      RECT 2.295 0.582 2.345 0.66 ;
      RECT 2.255 0.532 2.345 0.582 ;
    LAYER PO ;
      RECT 1.733 0.066 1.763 0.683 ;
      RECT 1.581 0.066 1.611 0.683 ;
      RECT 1.581 0.97 1.611 1.606 ;
      RECT 1.885 0.066 1.915 1.606 ;
      RECT 1.277 0.066 1.307 1.606 ;
      RECT 0.669 1.11 0.699 1.606 ;
      RECT 2.189 0.066 2.219 1.606 ;
      RECT 2.037 0.066 2.067 1.606 ;
      RECT 2.341 0.066 2.371 1.606 ;
      RECT 2.493 0.066 2.523 1.606 ;
      RECT 2.949 0.066 2.979 1.606 ;
      RECT 2.797 0.066 2.827 1.606 ;
      RECT 2.645 0.066 2.675 1.606 ;
      RECT 0.061 0.066 0.091 1.606 ;
      RECT 0.213 0.066 0.243 1.606 ;
      RECT 0.517 0.066 0.547 1.606 ;
      RECT 0.973 0.066 1.003 1.606 ;
      RECT 0.365 0.066 0.395 1.606 ;
      RECT 1.125 0.066 1.155 1.606 ;
      RECT 0.821 0.066 0.851 0.653 ;
      RECT 0.669 0.066 0.699 0.653 ;
      RECT 0.821 1.11 0.851 1.606 ;
      RECT 1.733 0.97 1.763 1.606 ;
      RECT 1.429 0.066 1.459 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 3.155 1.773 ;
  END
END DELLN1X2_RVT

MACRO DELLN2X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.952 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.679 0.401 0.721 ;
      LAYER M1 ;
        RECT 0.097 0.725 0.21 0.815 ;
        RECT 0.097 0.675 0.421 0.725 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0102 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.323 0.151 3.365 0.193 ;
        RECT 3.627 0.151 3.669 0.193 ;
        RECT 3.323 0.243 3.365 0.285 ;
        RECT 3.627 0.243 3.669 0.285 ;
        RECT 3.323 0.335 3.365 0.377 ;
        RECT 3.627 0.335 3.669 0.377 ;
        RECT 3.323 0.427 3.365 0.469 ;
        RECT 3.627 0.427 3.669 0.469 ;
        RECT 3.323 1.027 3.365 1.069 ;
        RECT 3.627 1.027 3.669 1.069 ;
        RECT 3.323 1.119 3.365 1.161 ;
        RECT 3.627 1.119 3.669 1.161 ;
        RECT 3.323 1.211 3.365 1.253 ;
        RECT 3.627 1.211 3.669 1.253 ;
        RECT 3.323 1.303 3.365 1.345 ;
        RECT 3.627 1.303 3.669 1.345 ;
        RECT 3.323 1.395 3.365 1.437 ;
        RECT 3.627 1.395 3.669 1.437 ;
        RECT 3.323 1.487 3.365 1.529 ;
        RECT 3.627 1.487 3.669 1.529 ;
      LAYER M1 ;
        RECT 3.319 0.942 3.369 1.564 ;
        RECT 3.623 0.942 3.673 1.564 ;
        RECT 3.319 0.892 3.729 0.942 ;
        RECT 3.679 0.663 3.729 0.892 ;
        RECT 3.679 0.587 3.855 0.663 ;
        RECT 3.319 0.537 3.855 0.587 ;
        RECT 3.319 0.116 3.369 0.537 ;
        RECT 3.623 0.116 3.673 0.537 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.663 0.603 0.705 0.645 ;
        RECT 0.815 0.603 0.857 0.645 ;
        RECT 1.575 0.603 1.617 0.645 ;
        RECT 1.727 0.603 1.769 0.645 ;
        RECT 2.487 0.603 2.529 0.645 ;
        RECT 2.639 0.603 2.681 0.645 ;
        RECT 2.107 0.81 2.149 0.852 ;
        RECT 0.283 0.827 0.325 0.869 ;
        RECT 3.019 0.836 3.061 0.878 ;
        RECT 1.195 0.837 1.237 0.879 ;
        RECT 2.107 0.902 2.149 0.944 ;
        RECT 2.411 0.906 2.453 0.948 ;
        RECT 0.283 0.919 0.325 0.961 ;
        RECT 3.019 0.928 3.061 0.97 ;
        RECT 1.195 0.929 1.237 0.971 ;
        RECT 2.411 0.998 2.453 1.04 ;
        RECT 3.019 1.02 3.061 1.062 ;
        RECT 3.475 1.027 3.517 1.069 ;
        RECT 2.411 1.09 2.453 1.132 ;
        RECT 3.019 1.112 3.061 1.154 ;
        RECT 3.475 1.119 3.517 1.161 ;
        RECT 2.411 1.182 2.453 1.224 ;
        RECT 0.587 1.2 0.629 1.242 ;
        RECT 3.019 1.204 3.061 1.246 ;
        RECT 3.475 1.211 3.517 1.253 ;
        RECT 2.411 1.274 2.453 1.316 ;
        RECT 0.587 1.292 0.629 1.334 ;
        RECT 1.499 1.3 1.541 1.342 ;
        RECT 3.475 1.303 3.517 1.345 ;
        RECT 2.411 1.366 2.453 1.408 ;
        RECT 0.587 1.384 0.629 1.426 ;
        RECT 1.499 1.392 1.541 1.434 ;
        RECT 3.475 1.395 3.517 1.437 ;
        RECT 0.587 1.476 0.629 1.518 ;
        RECT 1.499 1.484 1.541 1.526 ;
        RECT 3.475 1.487 3.517 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
        RECT 3.095 1.651 3.137 1.693 ;
        RECT 3.247 1.651 3.289 1.693 ;
        RECT 3.399 1.651 3.441 1.693 ;
        RECT 3.551 1.651 3.593 1.693 ;
        RECT 3.703 1.651 3.745 1.693 ;
        RECT 3.855 1.651 3.897 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 3.952 1.702 ;
        RECT 2.367 1.428 2.417 1.642 ;
        RECT 2.367 1.378 2.457 1.428 ;
        RECT 1.495 1.29 1.545 1.642 ;
        RECT 1.455 1.24 1.545 1.29 ;
        RECT 0.583 1.21 0.633 1.642 ;
        RECT 0.543 1.16 0.633 1.21 ;
        RECT 1.455 1.091 1.505 1.24 ;
        RECT 1.455 1.041 1.545 1.091 ;
        RECT 3.471 0.992 3.521 1.642 ;
        RECT 0.543 1.01 0.593 1.16 ;
        RECT 0.279 0.807 0.329 1.642 ;
        RECT 1.191 0.817 1.241 1.642 ;
        RECT 2.103 0.775 2.153 1.642 ;
        RECT 3.015 0.816 3.065 1.642 ;
        RECT 0.543 0.96 0.637 1.01 ;
        RECT 2.407 0.649 2.457 1.378 ;
        RECT 1.495 0.649 1.545 1.041 ;
        RECT 0.587 0.649 0.637 0.96 ;
        RECT 0.587 0.599 0.877 0.649 ;
        RECT 1.495 0.599 1.789 0.649 ;
        RECT 2.407 0.599 2.701 0.649 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 3.399 -0.021 3.441 0.021 ;
        RECT 3.551 -0.021 3.593 0.021 ;
        RECT 3.703 -0.021 3.745 0.021 ;
        RECT 3.855 -0.021 3.897 0.021 ;
        RECT 3.475 0.149 3.517 0.191 ;
        RECT 3.475 0.241 3.517 0.283 ;
        RECT 3.019 0.301 3.061 0.343 ;
        RECT 2.411 0.331 2.453 0.373 ;
        RECT 3.475 0.333 3.517 0.375 ;
        RECT 0.587 0.381 0.629 0.423 ;
        RECT 3.019 0.393 3.061 0.435 ;
        RECT 1.499 0.401 1.541 0.443 ;
        RECT 2.411 0.424 2.453 0.466 ;
        RECT 0.587 0.474 0.629 0.516 ;
        RECT 0.283 0.478 0.325 0.52 ;
        RECT 1.195 0.478 1.237 0.52 ;
        RECT 3.019 0.485 3.061 0.527 ;
        RECT 2.107 0.514 2.149 0.556 ;
        RECT 0.663 1.064 0.705 1.106 ;
        RECT 0.815 1.064 0.857 1.106 ;
        RECT 1.575 1.144 1.617 1.186 ;
        RECT 1.727 1.144 1.769 1.186 ;
        RECT 2.487 1.526 2.529 1.568 ;
        RECT 2.639 1.526 2.681 1.568 ;
      LAYER M1 ;
        RECT 2.467 1.522 2.801 1.572 ;
        RECT 1.555 1.14 1.889 1.19 ;
        RECT 0.643 1.06 0.977 1.11 ;
        RECT 2.751 0.549 2.801 1.522 ;
        RECT 1.839 0.549 1.889 1.14 ;
        RECT 0.927 0.549 0.977 1.06 ;
        RECT 0.583 0.499 0.977 0.549 ;
        RECT 1.495 0.499 1.889 0.549 ;
        RECT 2.407 0.499 2.801 0.549 ;
        RECT 2.103 0.316 2.153 0.58 ;
        RECT 2.103 0.266 2.156 0.316 ;
        RECT 0.583 0.248 0.633 0.499 ;
        RECT 1.495 0.248 1.545 0.499 ;
        RECT 2.407 0.248 2.457 0.499 ;
        RECT 0.583 0.198 1.129 0.248 ;
        RECT 1.495 0.198 2.041 0.248 ;
        RECT 2.407 0.198 2.953 0.248 ;
        RECT 3.015 0.03 3.065 0.547 ;
        RECT 0.279 0.03 0.329 0.54 ;
        RECT 1.191 0.03 1.241 0.54 ;
        RECT 3.471 0.03 3.521 0.41 ;
        RECT 2.106 0.03 2.156 0.266 ;
        RECT 1.079 0.03 1.129 0.198 ;
        RECT 1.991 0.03 2.041 0.198 ;
        RECT 2.903 0.03 2.953 0.198 ;
        RECT 0 -0.03 3.952 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 2.259 0.514 2.301 0.556 ;
      RECT 2.791 0.1 2.833 0.142 ;
      RECT 2.867 0.489 2.909 0.531 ;
      RECT 2.867 0.489 2.909 0.531 ;
      RECT 2.183 0.675 2.225 0.717 ;
      RECT 2.259 0.81 2.301 0.852 ;
      RECT 2.259 0.81 2.301 0.852 ;
      RECT 1.043 0.397 1.085 0.439 ;
      RECT 1.955 1.339 1.997 1.381 ;
      RECT 2.867 1.091 2.909 1.133 ;
      RECT 2.867 1.091 2.909 1.133 ;
      RECT 2.867 0.998 2.909 1.04 ;
      RECT 2.867 0.906 2.909 0.948 ;
      RECT 2.867 0.906 2.909 0.948 ;
      RECT 2.867 0.998 2.909 1.04 ;
      RECT 1.955 0.428 1.997 0.47 ;
      RECT 0.435 0.902 0.477 0.944 ;
      RECT 1.347 0.929 1.389 0.971 ;
      RECT 3.171 0.305 3.213 0.347 ;
      RECT 1.347 0.929 1.389 0.971 ;
      RECT 3.095 0.664 3.137 0.706 ;
      RECT 1.955 1.246 1.997 1.288 ;
      RECT 3.171 0.928 3.213 0.97 ;
      RECT 3.171 1.204 3.213 1.246 ;
      RECT 3.399 0.664 3.441 0.706 ;
      RECT 3.171 1.112 3.213 1.154 ;
      RECT 3.171 1.02 3.213 1.062 ;
      RECT 3.171 0.928 3.213 0.97 ;
      RECT 3.171 0.489 3.213 0.531 ;
      RECT 3.171 0.397 3.213 0.439 ;
      RECT 3.171 0.397 3.213 0.439 ;
      RECT 2.867 1.368 2.909 1.41 ;
      RECT 2.867 0.397 2.909 0.439 ;
      RECT 2.867 0.397 2.909 0.439 ;
      RECT 2.867 1.183 2.909 1.225 ;
      RECT 0.435 0.902 0.477 0.944 ;
      RECT 2.867 1.183 2.909 1.225 ;
      RECT 0.435 0.81 0.477 0.852 ;
      RECT 1.043 1.258 1.085 1.3 ;
      RECT 0.435 0.478 0.477 0.52 ;
      RECT 1.043 0.489 1.085 0.531 ;
      RECT 1.043 1.166 1.085 1.208 ;
      RECT 1.043 1.443 1.085 1.485 ;
      RECT 1.043 1.166 1.085 1.208 ;
      RECT 1.043 1.258 1.085 1.3 ;
      RECT 2.867 1.275 2.909 1.317 ;
      RECT 0.435 0.478 0.477 0.52 ;
      RECT 0.967 0.1 1.009 0.142 ;
      RECT 1.955 1.246 1.997 1.288 ;
      RECT 1.955 1.339 1.997 1.381 ;
      RECT 1.043 1.351 1.085 1.393 ;
      RECT 1.043 1.351 1.085 1.393 ;
      RECT 1.347 0.837 1.389 0.879 ;
      RECT 1.347 0.837 1.389 0.879 ;
      RECT 1.347 0.478 1.389 0.52 ;
      RECT 1.271 0.679 1.313 0.721 ;
      RECT 2.867 1.275 2.909 1.317 ;
      RECT 1.043 0.397 1.085 0.439 ;
      RECT 2.867 1.368 2.909 1.41 ;
      RECT 0.435 0.81 0.477 0.852 ;
      RECT 3.551 0.664 3.593 0.706 ;
      RECT 3.171 1.02 3.213 1.062 ;
      RECT 3.171 1.112 3.213 1.154 ;
      RECT 1.879 0.1 1.921 0.142 ;
      RECT 1.043 1.443 1.085 1.485 ;
      RECT 1.043 0.489 1.085 0.531 ;
      RECT 1.955 1.431 1.997 1.473 ;
      RECT 1.955 1.431 1.997 1.473 ;
      RECT 3.171 1.204 3.213 1.246 ;
      RECT 1.955 0.428 1.997 0.47 ;
    LAYER M1 ;
      RECT 3.207 0.66 3.628 0.71 ;
      RECT 3.167 0.285 3.217 0.532 ;
      RECT 3.167 0.532 3.257 0.582 ;
      RECT 3.167 0.887 3.257 0.937 ;
      RECT 3.167 0.937 3.217 1.266 ;
      RECT 3.207 0.71 3.257 0.887 ;
      RECT 3.207 0.582 3.257 0.66 ;
      RECT 2.863 0.66 3.157 0.71 ;
      RECT 2.863 0.71 2.913 1.43 ;
      RECT 2.863 0.377 2.913 0.66 ;
      RECT 2.255 0.096 2.853 0.146 ;
      RECT 2.255 0.532 2.345 0.582 ;
      RECT 2.255 0.825 2.305 0.887 ;
      RECT 2.255 0.775 2.345 0.825 ;
      RECT 2.255 0.146 2.305 0.532 ;
      RECT 2.295 0.582 2.345 0.775 ;
      RECT 1.039 0.675 1.333 0.725 ;
      RECT 1.039 0.725 1.089 1.505 ;
      RECT 1.039 0.377 1.089 0.675 ;
      RECT 0.431 0.096 1.029 0.146 ;
      RECT 0.431 0.541 0.521 0.591 ;
      RECT 0.431 0.146 0.481 0.541 ;
      RECT 0.431 0.775 0.521 0.825 ;
      RECT 0.431 0.825 0.481 0.964 ;
      RECT 0.471 0.591 0.521 0.775 ;
      RECT 1.951 0.671 2.245 0.721 ;
      RECT 1.951 0.721 2.001 1.493 ;
      RECT 1.951 0.381 2.001 0.671 ;
      RECT 1.343 0.096 1.941 0.146 ;
      RECT 1.343 0.532 1.433 0.582 ;
      RECT 1.343 0.775 1.433 0.825 ;
      RECT 1.343 0.146 1.393 0.532 ;
      RECT 1.343 0.825 1.393 0.991 ;
      RECT 1.383 0.582 1.433 0.775 ;
    LAYER PO ;
      RECT 0.213 0.066 0.243 1.606 ;
      RECT 2.493 0.066 2.523 0.683 ;
      RECT 2.493 0.826 2.523 1.606 ;
      RECT 2.645 0.066 2.675 0.683 ;
      RECT 2.645 0.826 2.675 1.606 ;
      RECT 0.517 0.066 0.547 1.606 ;
      RECT 0.973 0.066 1.003 1.606 ;
      RECT 0.365 0.066 0.395 1.606 ;
      RECT 1.125 0.066 1.155 1.606 ;
      RECT 0.821 0.066 0.851 0.683 ;
      RECT 0.669 0.066 0.699 0.683 ;
      RECT 0.821 1.03 0.851 1.606 ;
      RECT 1.733 1.11 1.763 1.606 ;
      RECT 1.429 0.066 1.459 1.606 ;
      RECT 1.733 0.066 1.763 0.683 ;
      RECT 1.581 0.066 1.611 0.683 ;
      RECT 1.581 1.11 1.611 1.606 ;
      RECT 1.885 0.066 1.915 1.606 ;
      RECT 3.253 0.066 3.283 1.606 ;
      RECT 1.277 0.066 1.307 1.606 ;
      RECT 3.557 0.066 3.587 1.606 ;
      RECT 3.101 0.066 3.131 1.606 ;
      RECT 3.709 0.066 3.739 1.606 ;
      RECT 3.405 0.066 3.435 1.606 ;
      RECT 3.861 0.066 3.891 1.606 ;
      RECT 0.669 1.03 0.699 1.606 ;
      RECT 2.189 0.066 2.219 1.606 ;
      RECT 2.037 0.066 2.067 1.606 ;
      RECT 2.341 0.066 2.371 1.606 ;
      RECT 0.061 0.066 0.091 1.606 ;
      RECT 2.949 0.066 2.979 1.606 ;
      RECT 2.797 0.066 2.827 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 4.067 1.773 ;
  END
END DELLN2X2_RVT

MACRO NBUFFX16_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.648 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.664 0.401 0.706 ;
        RECT 0.511 0.664 0.553 0.706 ;
        RECT 0.663 0.664 0.705 0.706 ;
      LAYER M1 ;
        RECT 0.249 0.71 0.362 0.815 ;
        RECT 0.249 0.66 0.74 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1098 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.891 0.151 0.933 0.193 ;
        RECT 1.195 0.151 1.237 0.193 ;
        RECT 1.499 0.151 1.541 0.193 ;
        RECT 1.803 0.151 1.845 0.193 ;
        RECT 2.411 0.151 2.453 0.193 ;
        RECT 2.715 0.151 2.757 0.193 ;
        RECT 3.019 0.151 3.061 0.193 ;
        RECT 3.323 0.151 3.365 0.193 ;
        RECT 2.107 0.152 2.149 0.194 ;
        RECT 0.891 0.243 0.933 0.285 ;
        RECT 1.195 0.243 1.237 0.285 ;
        RECT 1.499 0.243 1.541 0.285 ;
        RECT 1.803 0.243 1.845 0.285 ;
        RECT 2.411 0.243 2.453 0.285 ;
        RECT 2.715 0.243 2.757 0.285 ;
        RECT 3.019 0.243 3.061 0.285 ;
        RECT 3.323 0.243 3.365 0.285 ;
        RECT 2.107 0.244 2.149 0.286 ;
        RECT 0.891 0.335 0.933 0.377 ;
        RECT 1.195 0.335 1.237 0.377 ;
        RECT 1.499 0.335 1.541 0.377 ;
        RECT 1.803 0.335 1.845 0.377 ;
        RECT 2.411 0.335 2.453 0.377 ;
        RECT 2.715 0.335 2.757 0.377 ;
        RECT 3.019 0.335 3.061 0.377 ;
        RECT 3.323 0.335 3.365 0.377 ;
        RECT 2.107 0.336 2.149 0.378 ;
        RECT 0.891 0.427 0.933 0.469 ;
        RECT 1.195 0.427 1.237 0.469 ;
        RECT 1.499 0.427 1.541 0.469 ;
        RECT 1.803 0.427 1.845 0.469 ;
        RECT 2.411 0.427 2.453 0.469 ;
        RECT 2.715 0.427 2.757 0.469 ;
        RECT 3.019 0.427 3.061 0.469 ;
        RECT 3.323 0.427 3.365 0.469 ;
        RECT 2.107 0.428 2.149 0.47 ;
        RECT 0.891 1.027 0.933 1.069 ;
        RECT 1.195 1.027 1.237 1.069 ;
        RECT 1.499 1.027 1.541 1.069 ;
        RECT 1.803 1.027 1.845 1.069 ;
        RECT 2.411 1.027 2.453 1.069 ;
        RECT 2.715 1.027 2.757 1.069 ;
        RECT 3.019 1.027 3.061 1.069 ;
        RECT 3.323 1.027 3.365 1.069 ;
        RECT 2.107 1.028 2.149 1.07 ;
        RECT 0.891 1.119 0.933 1.161 ;
        RECT 1.195 1.119 1.237 1.161 ;
        RECT 1.499 1.119 1.541 1.161 ;
        RECT 1.803 1.119 1.845 1.161 ;
        RECT 2.411 1.119 2.453 1.161 ;
        RECT 2.715 1.119 2.757 1.161 ;
        RECT 3.019 1.119 3.061 1.161 ;
        RECT 3.323 1.119 3.365 1.161 ;
        RECT 2.107 1.12 2.149 1.162 ;
        RECT 0.891 1.211 0.933 1.253 ;
        RECT 1.195 1.211 1.237 1.253 ;
        RECT 1.499 1.211 1.541 1.253 ;
        RECT 1.803 1.211 1.845 1.253 ;
        RECT 2.411 1.211 2.453 1.253 ;
        RECT 2.715 1.211 2.757 1.253 ;
        RECT 3.019 1.211 3.061 1.253 ;
        RECT 3.323 1.211 3.365 1.253 ;
        RECT 2.107 1.212 2.149 1.254 ;
        RECT 0.891 1.303 0.933 1.345 ;
        RECT 1.195 1.303 1.237 1.345 ;
        RECT 1.499 1.303 1.541 1.345 ;
        RECT 1.803 1.303 1.845 1.345 ;
        RECT 2.411 1.303 2.453 1.345 ;
        RECT 2.715 1.303 2.757 1.345 ;
        RECT 3.019 1.303 3.061 1.345 ;
        RECT 3.323 1.303 3.365 1.345 ;
        RECT 2.107 1.304 2.149 1.346 ;
        RECT 0.891 1.395 0.933 1.437 ;
        RECT 1.195 1.395 1.237 1.437 ;
        RECT 1.499 1.395 1.541 1.437 ;
        RECT 1.803 1.395 1.845 1.437 ;
        RECT 2.411 1.395 2.453 1.437 ;
        RECT 2.715 1.395 2.757 1.437 ;
        RECT 3.019 1.395 3.061 1.437 ;
        RECT 3.323 1.395 3.365 1.437 ;
        RECT 2.107 1.396 2.149 1.438 ;
        RECT 0.891 1.487 0.933 1.529 ;
        RECT 1.195 1.487 1.237 1.529 ;
        RECT 1.499 1.487 1.541 1.529 ;
        RECT 1.803 1.487 1.845 1.529 ;
        RECT 2.411 1.487 2.453 1.529 ;
        RECT 2.715 1.487 2.757 1.529 ;
        RECT 3.019 1.487 3.061 1.529 ;
        RECT 3.323 1.487 3.365 1.529 ;
        RECT 2.107 1.488 2.149 1.53 ;
      LAYER M1 ;
        RECT 2.103 0.942 2.153 1.565 ;
        RECT 0.887 0.942 0.937 1.564 ;
        RECT 1.191 0.942 1.241 1.564 ;
        RECT 1.495 0.942 1.545 1.564 ;
        RECT 1.799 0.942 1.849 1.564 ;
        RECT 2.407 0.942 2.457 1.564 ;
        RECT 2.711 0.942 2.761 1.564 ;
        RECT 3.015 0.942 3.065 1.564 ;
        RECT 3.319 0.942 3.369 1.564 ;
        RECT 0.887 0.892 3.428 0.942 ;
        RECT 3.378 0.663 3.428 0.892 ;
        RECT 3.378 0.587 3.551 0.663 ;
        RECT 0.887 0.537 3.551 0.587 ;
        RECT 0.887 0.116 0.937 0.537 ;
        RECT 1.191 0.116 1.241 0.537 ;
        RECT 1.495 0.116 1.545 0.537 ;
        RECT 1.799 0.116 1.849 0.537 ;
        RECT 2.103 0.117 2.153 0.537 ;
        RECT 2.407 0.116 2.457 0.537 ;
        RECT 2.711 0.116 2.761 0.537 ;
        RECT 3.015 0.116 3.065 0.537 ;
        RECT 3.319 0.116 3.369 0.537 ;
    END
    ANTENNADIFFAREA 1.2904 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.435 1.027 0.477 1.069 ;
        RECT 0.739 1.027 0.781 1.069 ;
        RECT 1.043 1.027 1.085 1.069 ;
        RECT 1.347 1.027 1.389 1.069 ;
        RECT 1.651 1.027 1.693 1.069 ;
        RECT 1.955 1.027 1.997 1.069 ;
        RECT 2.259 1.027 2.301 1.069 ;
        RECT 2.563 1.027 2.605 1.069 ;
        RECT 2.867 1.027 2.909 1.069 ;
        RECT 3.171 1.027 3.213 1.069 ;
        RECT 0.435 1.119 0.477 1.161 ;
        RECT 0.739 1.119 0.781 1.161 ;
        RECT 1.043 1.119 1.085 1.161 ;
        RECT 1.347 1.119 1.389 1.161 ;
        RECT 1.651 1.119 1.693 1.161 ;
        RECT 1.955 1.119 1.997 1.161 ;
        RECT 2.259 1.119 2.301 1.161 ;
        RECT 2.563 1.119 2.605 1.161 ;
        RECT 2.867 1.119 2.909 1.161 ;
        RECT 3.171 1.119 3.213 1.161 ;
        RECT 0.435 1.211 0.477 1.253 ;
        RECT 0.739 1.211 0.781 1.253 ;
        RECT 1.043 1.211 1.085 1.253 ;
        RECT 1.347 1.211 1.389 1.253 ;
        RECT 1.651 1.211 1.693 1.253 ;
        RECT 1.955 1.211 1.997 1.253 ;
        RECT 2.259 1.211 2.301 1.253 ;
        RECT 2.563 1.211 2.605 1.253 ;
        RECT 2.867 1.211 2.909 1.253 ;
        RECT 3.171 1.211 3.213 1.253 ;
        RECT 0.435 1.303 0.477 1.345 ;
        RECT 0.739 1.303 0.781 1.345 ;
        RECT 1.043 1.303 1.085 1.345 ;
        RECT 1.347 1.303 1.389 1.345 ;
        RECT 1.651 1.303 1.693 1.345 ;
        RECT 1.955 1.303 1.997 1.345 ;
        RECT 2.259 1.303 2.301 1.345 ;
        RECT 2.563 1.303 2.605 1.345 ;
        RECT 2.867 1.303 2.909 1.345 ;
        RECT 3.171 1.303 3.213 1.345 ;
        RECT 0.435 1.395 0.477 1.437 ;
        RECT 0.739 1.395 0.781 1.437 ;
        RECT 1.043 1.395 1.085 1.437 ;
        RECT 1.347 1.395 1.389 1.437 ;
        RECT 1.651 1.395 1.693 1.437 ;
        RECT 1.955 1.395 1.997 1.437 ;
        RECT 2.259 1.395 2.301 1.437 ;
        RECT 2.563 1.395 2.605 1.437 ;
        RECT 2.867 1.395 2.909 1.437 ;
        RECT 3.171 1.395 3.213 1.437 ;
        RECT 0.435 1.487 0.477 1.529 ;
        RECT 0.739 1.487 0.781 1.529 ;
        RECT 1.043 1.487 1.085 1.529 ;
        RECT 1.347 1.487 1.389 1.529 ;
        RECT 1.651 1.487 1.693 1.529 ;
        RECT 1.955 1.487 1.997 1.529 ;
        RECT 2.259 1.487 2.301 1.529 ;
        RECT 2.563 1.487 2.605 1.529 ;
        RECT 2.867 1.487 2.909 1.529 ;
        RECT 3.171 1.487 3.213 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
        RECT 3.095 1.651 3.137 1.693 ;
        RECT 3.247 1.651 3.289 1.693 ;
        RECT 3.399 1.651 3.441 1.693 ;
        RECT 3.551 1.651 3.593 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 3.648 1.702 ;
        RECT 0.431 0.992 0.481 1.642 ;
        RECT 0.735 0.992 0.785 1.642 ;
        RECT 1.039 0.992 1.089 1.642 ;
        RECT 1.343 0.992 1.393 1.642 ;
        RECT 1.647 0.992 1.697 1.642 ;
        RECT 1.951 0.992 2.001 1.642 ;
        RECT 2.255 0.992 2.305 1.642 ;
        RECT 2.559 0.992 2.609 1.642 ;
        RECT 2.863 0.992 2.913 1.642 ;
        RECT 3.167 0.992 3.217 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 3.399 -0.021 3.441 0.021 ;
        RECT 3.551 -0.021 3.593 0.021 ;
        RECT 0.435 0.149 0.477 0.191 ;
        RECT 0.739 0.149 0.781 0.191 ;
        RECT 1.043 0.149 1.085 0.191 ;
        RECT 1.347 0.149 1.389 0.191 ;
        RECT 1.651 0.149 1.693 0.191 ;
        RECT 1.955 0.149 1.997 0.191 ;
        RECT 2.259 0.149 2.301 0.191 ;
        RECT 2.563 0.149 2.605 0.191 ;
        RECT 2.867 0.149 2.909 0.191 ;
        RECT 3.171 0.149 3.213 0.191 ;
        RECT 0.435 0.241 0.477 0.283 ;
        RECT 0.739 0.241 0.781 0.283 ;
        RECT 1.043 0.241 1.085 0.283 ;
        RECT 1.347 0.241 1.389 0.283 ;
        RECT 1.651 0.241 1.693 0.283 ;
        RECT 1.955 0.241 1.997 0.283 ;
        RECT 2.259 0.241 2.301 0.283 ;
        RECT 2.563 0.241 2.605 0.283 ;
        RECT 2.867 0.241 2.909 0.283 ;
        RECT 3.171 0.241 3.213 0.283 ;
        RECT 0.435 0.333 0.477 0.375 ;
        RECT 0.739 0.333 0.781 0.375 ;
        RECT 1.043 0.333 1.085 0.375 ;
        RECT 1.347 0.333 1.389 0.375 ;
        RECT 1.651 0.333 1.693 0.375 ;
        RECT 1.955 0.333 1.997 0.375 ;
        RECT 2.259 0.333 2.301 0.375 ;
        RECT 2.563 0.333 2.605 0.375 ;
        RECT 2.867 0.333 2.909 0.375 ;
        RECT 3.171 0.333 3.213 0.375 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.41 ;
        RECT 0.735 0.03 0.785 0.41 ;
        RECT 1.039 0.03 1.089 0.41 ;
        RECT 1.343 0.03 1.393 0.41 ;
        RECT 1.647 0.03 1.697 0.41 ;
        RECT 1.951 0.03 2.001 0.41 ;
        RECT 2.255 0.03 2.305 0.41 ;
        RECT 2.559 0.03 2.609 0.41 ;
        RECT 2.863 0.03 2.913 0.41 ;
        RECT 3.167 0.03 3.217 0.41 ;
        RECT 0 -0.03 3.648 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.587 0.151 0.629 0.193 ;
      RECT 0.587 1.027 0.629 1.069 ;
      RECT 0.587 0.427 0.629 0.469 ;
      RECT 0.587 0.335 0.629 0.377 ;
      RECT 0.587 1.119 0.629 1.161 ;
      RECT 0.587 1.027 0.629 1.069 ;
      RECT 0.587 0.335 0.629 0.377 ;
      RECT 0.587 1.487 0.629 1.529 ;
      RECT 0.587 0.243 0.629 0.285 ;
      RECT 0.587 1.487 0.629 1.529 ;
      RECT 0.587 1.395 0.629 1.437 ;
      RECT 0.587 0.151 0.629 0.193 ;
      RECT 0.587 1.119 0.629 1.161 ;
      RECT 0.587 1.395 0.629 1.437 ;
      RECT 0.587 1.211 0.629 1.253 ;
      RECT 0.587 1.211 0.629 1.253 ;
      RECT 0.587 1.303 0.629 1.345 ;
      RECT 0.587 1.303 0.629 1.345 ;
      RECT 0.283 1.027 0.325 1.069 ;
      RECT 0.283 1.119 0.325 1.161 ;
      RECT 0.283 1.027 0.325 1.069 ;
      RECT 0.283 1.487 0.325 1.529 ;
      RECT 0.283 1.487 0.325 1.529 ;
      RECT 0.283 1.395 0.325 1.437 ;
      RECT 0.283 1.119 0.325 1.161 ;
      RECT 0.283 1.395 0.325 1.437 ;
      RECT 0.283 1.211 0.325 1.253 ;
      RECT 0.283 1.211 0.325 1.253 ;
      RECT 0.283 1.303 0.325 1.345 ;
      RECT 0.283 1.303 0.325 1.345 ;
      RECT 0.283 0.151 0.325 0.193 ;
      RECT 0.283 0.427 0.325 0.469 ;
      RECT 0.283 0.335 0.325 0.377 ;
      RECT 0.283 0.335 0.325 0.377 ;
      RECT 0.283 0.243 0.325 0.285 ;
      RECT 0.283 0.151 0.325 0.193 ;
      RECT 2.183 0.664 2.225 0.706 ;
      RECT 2.639 0.664 2.681 0.706 ;
      RECT 2.335 0.664 2.377 0.706 ;
      RECT 2.487 0.664 2.529 0.706 ;
      RECT 2.031 0.664 2.073 0.706 ;
      RECT 2.791 0.664 2.833 0.706 ;
      RECT 3.247 0.664 3.289 0.706 ;
      RECT 2.943 0.664 2.985 0.706 ;
      RECT 3.095 0.664 3.137 0.706 ;
      RECT 1.727 0.664 1.769 0.706 ;
      RECT 1.879 0.664 1.921 0.706 ;
      RECT 1.575 0.664 1.617 0.706 ;
      RECT 1.423 0.664 1.465 0.706 ;
      RECT 1.271 0.664 1.313 0.706 ;
      RECT 0.967 0.664 1.009 0.706 ;
      RECT 1.119 0.664 1.161 0.706 ;
    LAYER M1 ;
      RECT 0.79 0.66 3.324 0.71 ;
      RECT 0.279 0.892 0.329 1.564 ;
      RECT 0.279 0.502 0.329 0.537 ;
      RECT 0.279 0.116 0.329 0.576 ;
      RECT 0.583 0.892 0.633 1.564 ;
      RECT 0.583 0.116 0.633 0.556 ;
      RECT 0.329 0.931 0.836 0.942 ;
      RECT 0.279 0.892 0.836 0.931 ;
      RECT 0.786 0.842 0.836 0.942 ;
      RECT 0.79 0.605 0.84 0.874 ;
      RECT 0.787 0.537 0.837 0.633 ;
      RECT 0.279 0.537 0.837 0.587 ;
    LAYER PO ;
      RECT 0.821 0.069 0.851 1.606 ;
      RECT 0.973 0.069 1.003 1.606 ;
      RECT 1.429 0.069 1.459 1.606 ;
      RECT 1.277 0.069 1.307 1.606 ;
      RECT 1.125 0.069 1.155 1.606 ;
      RECT 0.061 0.071 0.091 1.606 ;
      RECT 0.517 0.069 0.547 1.606 ;
      RECT 0.669 0.069 0.699 1.606 ;
      RECT 0.365 0.069 0.395 1.606 ;
      RECT 0.213 0.071 0.243 1.606 ;
      RECT 3.405 0.069 3.435 1.606 ;
      RECT 3.557 0.069 3.587 1.606 ;
      RECT 3.253 0.069 3.283 1.606 ;
      RECT 2.037 0.069 2.067 1.606 ;
      RECT 2.189 0.069 2.219 1.606 ;
      RECT 2.341 0.069 2.371 1.606 ;
      RECT 2.949 0.069 2.979 1.606 ;
      RECT 2.797 0.069 2.827 1.606 ;
      RECT 2.645 0.069 2.675 1.606 ;
      RECT 2.493 0.069 2.523 1.606 ;
      RECT 3.101 0.069 3.131 1.606 ;
      RECT 1.885 0.069 1.915 1.606 ;
      RECT 1.733 0.069 1.763 1.606 ;
      RECT 1.581 0.069 1.611 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 3.763 1.773 ;
  END
END NBUFFX16_RVT

MACRO NBUFFX32_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 6.384 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.664 0.401 0.706 ;
        RECT 0.511 0.664 0.553 0.706 ;
        RECT 0.663 0.664 0.705 0.706 ;
        RECT 0.815 0.664 0.857 0.706 ;
        RECT 0.967 0.664 1.009 0.706 ;
      LAYER M1 ;
        RECT 0.249 0.71 0.362 0.815 ;
        RECT 0.249 0.66 1.044 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.183 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.195 0.151 1.237 0.193 ;
        RECT 1.499 0.151 1.541 0.193 ;
        RECT 1.803 0.151 1.845 0.193 ;
        RECT 2.107 0.151 2.149 0.193 ;
        RECT 2.715 0.151 2.757 0.193 ;
        RECT 3.019 0.151 3.061 0.193 ;
        RECT 3.323 0.151 3.365 0.193 ;
        RECT 3.627 0.151 3.669 0.193 ;
        RECT 3.931 0.151 3.973 0.193 ;
        RECT 4.235 0.151 4.277 0.193 ;
        RECT 4.539 0.151 4.581 0.193 ;
        RECT 4.843 0.151 4.885 0.193 ;
        RECT 5.147 0.151 5.189 0.193 ;
        RECT 5.451 0.151 5.493 0.193 ;
        RECT 5.755 0.151 5.797 0.193 ;
        RECT 6.059 0.151 6.101 0.193 ;
        RECT 2.411 0.152 2.453 0.194 ;
        RECT 1.195 0.243 1.237 0.285 ;
        RECT 1.499 0.243 1.541 0.285 ;
        RECT 1.803 0.243 1.845 0.285 ;
        RECT 2.107 0.243 2.149 0.285 ;
        RECT 2.715 0.243 2.757 0.285 ;
        RECT 3.019 0.243 3.061 0.285 ;
        RECT 3.323 0.243 3.365 0.285 ;
        RECT 3.627 0.243 3.669 0.285 ;
        RECT 3.931 0.243 3.973 0.285 ;
        RECT 4.235 0.243 4.277 0.285 ;
        RECT 4.539 0.243 4.581 0.285 ;
        RECT 4.843 0.243 4.885 0.285 ;
        RECT 5.147 0.243 5.189 0.285 ;
        RECT 5.451 0.243 5.493 0.285 ;
        RECT 5.755 0.243 5.797 0.285 ;
        RECT 6.059 0.243 6.101 0.285 ;
        RECT 2.411 0.244 2.453 0.286 ;
        RECT 1.195 0.335 1.237 0.377 ;
        RECT 1.499 0.335 1.541 0.377 ;
        RECT 1.803 0.335 1.845 0.377 ;
        RECT 2.107 0.335 2.149 0.377 ;
        RECT 2.715 0.335 2.757 0.377 ;
        RECT 3.019 0.335 3.061 0.377 ;
        RECT 3.323 0.335 3.365 0.377 ;
        RECT 3.627 0.335 3.669 0.377 ;
        RECT 3.931 0.335 3.973 0.377 ;
        RECT 4.235 0.335 4.277 0.377 ;
        RECT 4.539 0.335 4.581 0.377 ;
        RECT 4.843 0.335 4.885 0.377 ;
        RECT 5.147 0.335 5.189 0.377 ;
        RECT 5.451 0.335 5.493 0.377 ;
        RECT 5.755 0.335 5.797 0.377 ;
        RECT 6.059 0.335 6.101 0.377 ;
        RECT 2.411 0.336 2.453 0.378 ;
        RECT 1.195 0.427 1.237 0.469 ;
        RECT 1.499 0.427 1.541 0.469 ;
        RECT 1.803 0.427 1.845 0.469 ;
        RECT 2.107 0.427 2.149 0.469 ;
        RECT 2.715 0.427 2.757 0.469 ;
        RECT 3.019 0.427 3.061 0.469 ;
        RECT 3.323 0.427 3.365 0.469 ;
        RECT 3.627 0.427 3.669 0.469 ;
        RECT 3.931 0.427 3.973 0.469 ;
        RECT 4.235 0.427 4.277 0.469 ;
        RECT 4.539 0.427 4.581 0.469 ;
        RECT 4.843 0.427 4.885 0.469 ;
        RECT 5.147 0.427 5.189 0.469 ;
        RECT 5.451 0.427 5.493 0.469 ;
        RECT 5.755 0.427 5.797 0.469 ;
        RECT 6.059 0.427 6.101 0.469 ;
        RECT 2.411 0.428 2.453 0.47 ;
        RECT 1.195 1.027 1.237 1.069 ;
        RECT 1.499 1.027 1.541 1.069 ;
        RECT 1.803 1.027 1.845 1.069 ;
        RECT 2.107 1.027 2.149 1.069 ;
        RECT 2.715 1.027 2.757 1.069 ;
        RECT 3.019 1.027 3.061 1.069 ;
        RECT 3.323 1.027 3.365 1.069 ;
        RECT 3.627 1.027 3.669 1.069 ;
        RECT 3.931 1.027 3.973 1.069 ;
        RECT 4.235 1.027 4.277 1.069 ;
        RECT 4.539 1.027 4.581 1.069 ;
        RECT 4.843 1.027 4.885 1.069 ;
        RECT 5.147 1.027 5.189 1.069 ;
        RECT 5.451 1.027 5.493 1.069 ;
        RECT 5.755 1.027 5.797 1.069 ;
        RECT 6.059 1.027 6.101 1.069 ;
        RECT 2.411 1.028 2.453 1.07 ;
        RECT 1.195 1.119 1.237 1.161 ;
        RECT 1.499 1.119 1.541 1.161 ;
        RECT 1.803 1.119 1.845 1.161 ;
        RECT 2.107 1.119 2.149 1.161 ;
        RECT 2.715 1.119 2.757 1.161 ;
        RECT 3.019 1.119 3.061 1.161 ;
        RECT 3.323 1.119 3.365 1.161 ;
        RECT 3.627 1.119 3.669 1.161 ;
        RECT 3.931 1.119 3.973 1.161 ;
        RECT 4.235 1.119 4.277 1.161 ;
        RECT 4.539 1.119 4.581 1.161 ;
        RECT 4.843 1.119 4.885 1.161 ;
        RECT 5.147 1.119 5.189 1.161 ;
        RECT 5.451 1.119 5.493 1.161 ;
        RECT 5.755 1.119 5.797 1.161 ;
        RECT 6.059 1.119 6.101 1.161 ;
        RECT 2.411 1.12 2.453 1.162 ;
        RECT 1.195 1.211 1.237 1.253 ;
        RECT 1.499 1.211 1.541 1.253 ;
        RECT 1.803 1.211 1.845 1.253 ;
        RECT 2.107 1.211 2.149 1.253 ;
        RECT 2.715 1.211 2.757 1.253 ;
        RECT 3.019 1.211 3.061 1.253 ;
        RECT 3.323 1.211 3.365 1.253 ;
        RECT 3.627 1.211 3.669 1.253 ;
        RECT 3.931 1.211 3.973 1.253 ;
        RECT 4.235 1.211 4.277 1.253 ;
        RECT 4.539 1.211 4.581 1.253 ;
        RECT 4.843 1.211 4.885 1.253 ;
        RECT 5.147 1.211 5.189 1.253 ;
        RECT 5.451 1.211 5.493 1.253 ;
        RECT 5.755 1.211 5.797 1.253 ;
        RECT 6.059 1.211 6.101 1.253 ;
        RECT 2.411 1.212 2.453 1.254 ;
        RECT 1.195 1.303 1.237 1.345 ;
        RECT 1.499 1.303 1.541 1.345 ;
        RECT 1.803 1.303 1.845 1.345 ;
        RECT 2.107 1.303 2.149 1.345 ;
        RECT 2.715 1.303 2.757 1.345 ;
        RECT 3.019 1.303 3.061 1.345 ;
        RECT 3.323 1.303 3.365 1.345 ;
        RECT 3.627 1.303 3.669 1.345 ;
        RECT 3.931 1.303 3.973 1.345 ;
        RECT 4.235 1.303 4.277 1.345 ;
        RECT 4.539 1.303 4.581 1.345 ;
        RECT 4.843 1.303 4.885 1.345 ;
        RECT 5.147 1.303 5.189 1.345 ;
        RECT 5.451 1.303 5.493 1.345 ;
        RECT 5.755 1.303 5.797 1.345 ;
        RECT 6.059 1.303 6.101 1.345 ;
        RECT 2.411 1.304 2.453 1.346 ;
        RECT 1.195 1.395 1.237 1.437 ;
        RECT 1.499 1.395 1.541 1.437 ;
        RECT 1.803 1.395 1.845 1.437 ;
        RECT 2.107 1.395 2.149 1.437 ;
        RECT 2.715 1.395 2.757 1.437 ;
        RECT 3.019 1.395 3.061 1.437 ;
        RECT 3.323 1.395 3.365 1.437 ;
        RECT 3.627 1.395 3.669 1.437 ;
        RECT 3.931 1.395 3.973 1.437 ;
        RECT 4.235 1.395 4.277 1.437 ;
        RECT 4.539 1.395 4.581 1.437 ;
        RECT 4.843 1.395 4.885 1.437 ;
        RECT 5.147 1.395 5.189 1.437 ;
        RECT 5.451 1.395 5.493 1.437 ;
        RECT 5.755 1.395 5.797 1.437 ;
        RECT 6.059 1.395 6.101 1.437 ;
        RECT 2.411 1.396 2.453 1.438 ;
        RECT 1.195 1.487 1.237 1.529 ;
        RECT 1.499 1.487 1.541 1.529 ;
        RECT 1.803 1.487 1.845 1.529 ;
        RECT 2.107 1.487 2.149 1.529 ;
        RECT 2.715 1.487 2.757 1.529 ;
        RECT 3.019 1.487 3.061 1.529 ;
        RECT 3.323 1.487 3.365 1.529 ;
        RECT 3.627 1.487 3.669 1.529 ;
        RECT 3.931 1.487 3.973 1.529 ;
        RECT 4.235 1.487 4.277 1.529 ;
        RECT 4.539 1.487 4.581 1.529 ;
        RECT 4.843 1.487 4.885 1.529 ;
        RECT 5.147 1.487 5.189 1.529 ;
        RECT 5.451 1.487 5.493 1.529 ;
        RECT 5.755 1.487 5.797 1.529 ;
        RECT 6.059 1.487 6.101 1.529 ;
        RECT 2.411 1.488 2.453 1.53 ;
      LAYER M1 ;
        RECT 3.927 0.942 3.977 1.564 ;
        RECT 4.231 0.942 4.281 1.564 ;
        RECT 4.535 0.942 4.585 1.564 ;
        RECT 4.839 0.942 4.889 1.564 ;
        RECT 5.143 0.942 5.193 1.564 ;
        RECT 5.447 0.942 5.497 1.564 ;
        RECT 5.751 0.942 5.801 1.564 ;
        RECT 6.055 0.942 6.105 1.564 ;
        RECT 6.114 0.663 6.164 0.892 ;
        RECT 1.191 0.892 6.164 0.942 ;
        RECT 2.407 0.942 2.457 1.565 ;
        RECT 1.191 0.942 1.241 1.564 ;
        RECT 1.495 0.942 1.545 1.564 ;
        RECT 1.799 0.942 1.849 1.564 ;
        RECT 2.103 0.942 2.153 1.564 ;
        RECT 2.711 0.942 2.761 1.564 ;
        RECT 3.015 0.942 3.065 1.564 ;
        RECT 3.319 0.942 3.369 1.564 ;
        RECT 3.623 0.942 3.673 1.564 ;
        RECT 6.114 0.587 6.287 0.663 ;
        RECT 1.191 0.537 6.287 0.587 ;
        RECT 3.927 0.116 3.977 0.537 ;
        RECT 4.231 0.116 4.281 0.537 ;
        RECT 4.535 0.116 4.585 0.537 ;
        RECT 4.839 0.116 4.889 0.537 ;
        RECT 5.143 0.116 5.193 0.537 ;
        RECT 5.447 0.116 5.497 0.537 ;
        RECT 5.751 0.116 5.801 0.537 ;
        RECT 6.055 0.116 6.105 0.537 ;
        RECT 1.191 0.116 1.241 0.537 ;
        RECT 1.495 0.116 1.545 0.537 ;
        RECT 1.799 0.116 1.849 0.537 ;
        RECT 2.103 0.116 2.153 0.537 ;
        RECT 2.407 0.117 2.457 0.537 ;
        RECT 2.711 0.116 2.761 0.537 ;
        RECT 3.015 0.116 3.065 0.537 ;
        RECT 3.319 0.116 3.369 0.537 ;
        RECT 3.623 0.116 3.673 0.537 ;
    END
    ANTENNADIFFAREA 2.4808 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.435 1.027 0.477 1.069 ;
        RECT 0.739 1.027 0.781 1.069 ;
        RECT 1.043 1.027 1.085 1.069 ;
        RECT 1.347 1.027 1.389 1.069 ;
        RECT 1.651 1.027 1.693 1.069 ;
        RECT 1.955 1.027 1.997 1.069 ;
        RECT 2.259 1.027 2.301 1.069 ;
        RECT 2.563 1.027 2.605 1.069 ;
        RECT 2.867 1.027 2.909 1.069 ;
        RECT 3.171 1.027 3.213 1.069 ;
        RECT 3.475 1.027 3.517 1.069 ;
        RECT 3.779 1.027 3.821 1.069 ;
        RECT 4.083 1.027 4.125 1.069 ;
        RECT 4.387 1.027 4.429 1.069 ;
        RECT 4.691 1.027 4.733 1.069 ;
        RECT 4.995 1.027 5.037 1.069 ;
        RECT 5.299 1.027 5.341 1.069 ;
        RECT 5.603 1.027 5.645 1.069 ;
        RECT 5.907 1.027 5.949 1.069 ;
        RECT 0.435 1.119 0.477 1.161 ;
        RECT 0.739 1.119 0.781 1.161 ;
        RECT 1.043 1.119 1.085 1.161 ;
        RECT 1.347 1.119 1.389 1.161 ;
        RECT 1.651 1.119 1.693 1.161 ;
        RECT 1.955 1.119 1.997 1.161 ;
        RECT 2.259 1.119 2.301 1.161 ;
        RECT 2.563 1.119 2.605 1.161 ;
        RECT 2.867 1.119 2.909 1.161 ;
        RECT 3.171 1.119 3.213 1.161 ;
        RECT 3.475 1.119 3.517 1.161 ;
        RECT 3.779 1.119 3.821 1.161 ;
        RECT 4.083 1.119 4.125 1.161 ;
        RECT 4.387 1.119 4.429 1.161 ;
        RECT 4.691 1.119 4.733 1.161 ;
        RECT 4.995 1.119 5.037 1.161 ;
        RECT 5.299 1.119 5.341 1.161 ;
        RECT 5.603 1.119 5.645 1.161 ;
        RECT 5.907 1.119 5.949 1.161 ;
        RECT 0.435 1.211 0.477 1.253 ;
        RECT 0.739 1.211 0.781 1.253 ;
        RECT 1.043 1.211 1.085 1.253 ;
        RECT 1.347 1.211 1.389 1.253 ;
        RECT 1.651 1.211 1.693 1.253 ;
        RECT 1.955 1.211 1.997 1.253 ;
        RECT 2.259 1.211 2.301 1.253 ;
        RECT 2.563 1.211 2.605 1.253 ;
        RECT 2.867 1.211 2.909 1.253 ;
        RECT 3.171 1.211 3.213 1.253 ;
        RECT 3.475 1.211 3.517 1.253 ;
        RECT 3.779 1.211 3.821 1.253 ;
        RECT 4.083 1.211 4.125 1.253 ;
        RECT 4.387 1.211 4.429 1.253 ;
        RECT 4.691 1.211 4.733 1.253 ;
        RECT 4.995 1.211 5.037 1.253 ;
        RECT 5.299 1.211 5.341 1.253 ;
        RECT 5.603 1.211 5.645 1.253 ;
        RECT 5.907 1.211 5.949 1.253 ;
        RECT 0.435 1.303 0.477 1.345 ;
        RECT 0.739 1.303 0.781 1.345 ;
        RECT 1.043 1.303 1.085 1.345 ;
        RECT 1.347 1.303 1.389 1.345 ;
        RECT 1.651 1.303 1.693 1.345 ;
        RECT 1.955 1.303 1.997 1.345 ;
        RECT 2.259 1.303 2.301 1.345 ;
        RECT 2.563 1.303 2.605 1.345 ;
        RECT 2.867 1.303 2.909 1.345 ;
        RECT 3.171 1.303 3.213 1.345 ;
        RECT 3.475 1.303 3.517 1.345 ;
        RECT 3.779 1.303 3.821 1.345 ;
        RECT 4.083 1.303 4.125 1.345 ;
        RECT 4.387 1.303 4.429 1.345 ;
        RECT 4.691 1.303 4.733 1.345 ;
        RECT 4.995 1.303 5.037 1.345 ;
        RECT 5.299 1.303 5.341 1.345 ;
        RECT 5.603 1.303 5.645 1.345 ;
        RECT 5.907 1.303 5.949 1.345 ;
        RECT 0.435 1.395 0.477 1.437 ;
        RECT 0.739 1.395 0.781 1.437 ;
        RECT 1.043 1.395 1.085 1.437 ;
        RECT 1.347 1.395 1.389 1.437 ;
        RECT 1.651 1.395 1.693 1.437 ;
        RECT 1.955 1.395 1.997 1.437 ;
        RECT 2.259 1.395 2.301 1.437 ;
        RECT 2.563 1.395 2.605 1.437 ;
        RECT 2.867 1.395 2.909 1.437 ;
        RECT 3.171 1.395 3.213 1.437 ;
        RECT 3.475 1.395 3.517 1.437 ;
        RECT 3.779 1.395 3.821 1.437 ;
        RECT 4.083 1.395 4.125 1.437 ;
        RECT 4.387 1.395 4.429 1.437 ;
        RECT 4.691 1.395 4.733 1.437 ;
        RECT 4.995 1.395 5.037 1.437 ;
        RECT 5.299 1.395 5.341 1.437 ;
        RECT 5.603 1.395 5.645 1.437 ;
        RECT 5.907 1.395 5.949 1.437 ;
        RECT 0.435 1.487 0.477 1.529 ;
        RECT 0.739 1.487 0.781 1.529 ;
        RECT 1.043 1.487 1.085 1.529 ;
        RECT 1.347 1.487 1.389 1.529 ;
        RECT 1.651 1.487 1.693 1.529 ;
        RECT 1.955 1.487 1.997 1.529 ;
        RECT 2.259 1.487 2.301 1.529 ;
        RECT 2.563 1.487 2.605 1.529 ;
        RECT 2.867 1.487 2.909 1.529 ;
        RECT 3.171 1.487 3.213 1.529 ;
        RECT 3.475 1.487 3.517 1.529 ;
        RECT 3.779 1.487 3.821 1.529 ;
        RECT 4.083 1.487 4.125 1.529 ;
        RECT 4.387 1.487 4.429 1.529 ;
        RECT 4.691 1.487 4.733 1.529 ;
        RECT 4.995 1.487 5.037 1.529 ;
        RECT 5.299 1.487 5.341 1.529 ;
        RECT 5.603 1.487 5.645 1.529 ;
        RECT 5.907 1.487 5.949 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
        RECT 3.095 1.651 3.137 1.693 ;
        RECT 3.247 1.651 3.289 1.693 ;
        RECT 3.399 1.651 3.441 1.693 ;
        RECT 3.551 1.651 3.593 1.693 ;
        RECT 3.703 1.651 3.745 1.693 ;
        RECT 3.855 1.651 3.897 1.693 ;
        RECT 4.007 1.651 4.049 1.693 ;
        RECT 4.159 1.651 4.201 1.693 ;
        RECT 4.311 1.651 4.353 1.693 ;
        RECT 4.463 1.651 4.505 1.693 ;
        RECT 4.615 1.651 4.657 1.693 ;
        RECT 4.767 1.651 4.809 1.693 ;
        RECT 4.919 1.651 4.961 1.693 ;
        RECT 5.071 1.651 5.113 1.693 ;
        RECT 5.223 1.651 5.265 1.693 ;
        RECT 5.375 1.651 5.417 1.693 ;
        RECT 5.527 1.651 5.569 1.693 ;
        RECT 5.679 1.651 5.721 1.693 ;
        RECT 5.831 1.651 5.873 1.693 ;
        RECT 5.983 1.651 6.025 1.693 ;
        RECT 6.135 1.651 6.177 1.693 ;
        RECT 6.287 1.651 6.329 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 6.384 1.702 ;
        RECT 3.167 0.992 3.217 1.642 ;
        RECT 3.471 0.992 3.521 1.642 ;
        RECT 3.775 0.992 3.825 1.642 ;
        RECT 4.079 0.992 4.129 1.642 ;
        RECT 4.383 0.992 4.433 1.642 ;
        RECT 4.687 0.992 4.737 1.642 ;
        RECT 4.991 0.992 5.041 1.642 ;
        RECT 5.295 0.992 5.345 1.642 ;
        RECT 5.599 0.992 5.649 1.642 ;
        RECT 5.903 0.992 5.953 1.642 ;
        RECT 0.431 0.992 0.481 1.642 ;
        RECT 0.735 0.992 0.785 1.642 ;
        RECT 1.039 0.992 1.089 1.642 ;
        RECT 1.343 0.992 1.393 1.642 ;
        RECT 1.647 0.992 1.697 1.642 ;
        RECT 1.951 0.992 2.001 1.642 ;
        RECT 2.255 0.992 2.305 1.642 ;
        RECT 2.559 0.992 2.609 1.642 ;
        RECT 2.863 0.992 2.913 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 3.399 -0.021 3.441 0.021 ;
        RECT 3.551 -0.021 3.593 0.021 ;
        RECT 3.703 -0.021 3.745 0.021 ;
        RECT 3.855 -0.021 3.897 0.021 ;
        RECT 4.007 -0.021 4.049 0.021 ;
        RECT 4.159 -0.021 4.201 0.021 ;
        RECT 4.311 -0.021 4.353 0.021 ;
        RECT 4.463 -0.021 4.505 0.021 ;
        RECT 4.615 -0.021 4.657 0.021 ;
        RECT 4.767 -0.021 4.809 0.021 ;
        RECT 4.919 -0.021 4.961 0.021 ;
        RECT 5.071 -0.021 5.113 0.021 ;
        RECT 5.223 -0.021 5.265 0.021 ;
        RECT 5.375 -0.021 5.417 0.021 ;
        RECT 5.527 -0.021 5.569 0.021 ;
        RECT 5.679 -0.021 5.721 0.021 ;
        RECT 5.831 -0.021 5.873 0.021 ;
        RECT 5.983 -0.021 6.025 0.021 ;
        RECT 6.135 -0.021 6.177 0.021 ;
        RECT 6.287 -0.021 6.329 0.021 ;
        RECT 0.435 0.149 0.477 0.191 ;
        RECT 0.739 0.149 0.781 0.191 ;
        RECT 1.043 0.149 1.085 0.191 ;
        RECT 1.347 0.149 1.389 0.191 ;
        RECT 1.651 0.149 1.693 0.191 ;
        RECT 1.955 0.149 1.997 0.191 ;
        RECT 2.259 0.149 2.301 0.191 ;
        RECT 2.563 0.149 2.605 0.191 ;
        RECT 2.867 0.149 2.909 0.191 ;
        RECT 3.171 0.149 3.213 0.191 ;
        RECT 3.475 0.149 3.517 0.191 ;
        RECT 3.779 0.149 3.821 0.191 ;
        RECT 4.083 0.149 4.125 0.191 ;
        RECT 4.387 0.149 4.429 0.191 ;
        RECT 4.691 0.149 4.733 0.191 ;
        RECT 4.995 0.149 5.037 0.191 ;
        RECT 5.299 0.149 5.341 0.191 ;
        RECT 5.603 0.149 5.645 0.191 ;
        RECT 5.907 0.149 5.949 0.191 ;
        RECT 0.435 0.241 0.477 0.283 ;
        RECT 0.739 0.241 0.781 0.283 ;
        RECT 1.043 0.241 1.085 0.283 ;
        RECT 1.347 0.241 1.389 0.283 ;
        RECT 1.651 0.241 1.693 0.283 ;
        RECT 1.955 0.241 1.997 0.283 ;
        RECT 2.259 0.241 2.301 0.283 ;
        RECT 2.563 0.241 2.605 0.283 ;
        RECT 2.867 0.241 2.909 0.283 ;
        RECT 3.171 0.241 3.213 0.283 ;
        RECT 3.475 0.241 3.517 0.283 ;
        RECT 3.779 0.241 3.821 0.283 ;
        RECT 4.083 0.241 4.125 0.283 ;
        RECT 4.387 0.241 4.429 0.283 ;
        RECT 4.691 0.241 4.733 0.283 ;
        RECT 4.995 0.241 5.037 0.283 ;
        RECT 5.299 0.241 5.341 0.283 ;
        RECT 5.603 0.241 5.645 0.283 ;
        RECT 5.907 0.241 5.949 0.283 ;
        RECT 0.435 0.333 0.477 0.375 ;
        RECT 0.739 0.333 0.781 0.375 ;
        RECT 1.043 0.333 1.085 0.375 ;
        RECT 1.347 0.333 1.389 0.375 ;
        RECT 1.651 0.333 1.693 0.375 ;
        RECT 1.955 0.333 1.997 0.375 ;
        RECT 2.259 0.333 2.301 0.375 ;
        RECT 2.563 0.333 2.605 0.375 ;
        RECT 2.867 0.333 2.909 0.375 ;
        RECT 3.171 0.333 3.213 0.375 ;
        RECT 3.475 0.333 3.517 0.375 ;
        RECT 3.779 0.333 3.821 0.375 ;
        RECT 4.083 0.333 4.125 0.375 ;
        RECT 4.387 0.333 4.429 0.375 ;
        RECT 4.691 0.333 4.733 0.375 ;
        RECT 4.995 0.333 5.037 0.375 ;
        RECT 5.299 0.333 5.341 0.375 ;
        RECT 5.603 0.333 5.645 0.375 ;
        RECT 5.907 0.333 5.949 0.375 ;
      LAYER M1 ;
        RECT 3.167 0.03 3.217 0.41 ;
        RECT 0 -0.03 6.384 0.03 ;
        RECT 3.471 0.03 3.521 0.41 ;
        RECT 3.775 0.03 3.825 0.41 ;
        RECT 4.079 0.03 4.129 0.41 ;
        RECT 4.383 0.03 4.433 0.41 ;
        RECT 4.687 0.03 4.737 0.41 ;
        RECT 4.991 0.03 5.041 0.41 ;
        RECT 5.295 0.03 5.345 0.41 ;
        RECT 5.599 0.03 5.649 0.41 ;
        RECT 5.903 0.03 5.953 0.41 ;
        RECT 0.431 0.03 0.481 0.41 ;
        RECT 0.735 0.03 0.785 0.41 ;
        RECT 1.039 0.03 1.089 0.41 ;
        RECT 1.343 0.03 1.393 0.41 ;
        RECT 1.647 0.03 1.697 0.41 ;
        RECT 1.951 0.03 2.001 0.41 ;
        RECT 2.255 0.03 2.305 0.41 ;
        RECT 2.559 0.03 2.609 0.41 ;
        RECT 2.863 0.03 2.913 0.41 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.094 0.66 6.06 0.71 ;
      RECT 0.279 0.892 0.329 1.564 ;
      RECT 0.279 0.502 0.329 0.537 ;
      RECT 0.279 0.116 0.329 0.576 ;
      RECT 0.583 0.892 0.633 1.564 ;
      RECT 0.583 0.116 0.633 0.576 ;
      RECT 0.887 0.892 0.937 1.564 ;
      RECT 0.887 0.116 0.937 0.576 ;
      RECT 0.329 0.931 1.141 0.942 ;
      RECT 0.279 0.892 1.141 0.931 ;
      RECT 1.091 0.818 1.141 0.942 ;
      RECT 1.094 0.605 1.144 0.874 ;
      RECT 1.091 0.538 1.141 0.631 ;
      RECT 0.279 0.537 1.141 0.587 ;
    LAYER CO ;
      RECT 5.983 0.664 6.025 0.706 ;
      RECT 4.615 0.664 4.657 0.706 ;
      RECT 4.311 0.664 4.353 0.706 ;
      RECT 4.463 0.664 4.505 0.706 ;
      RECT 4.159 0.664 4.201 0.706 ;
      RECT 4.007 0.664 4.049 0.706 ;
      RECT 3.855 0.664 3.897 0.706 ;
      RECT 3.703 0.664 3.745 0.706 ;
      RECT 5.375 0.664 5.417 0.706 ;
      RECT 5.831 0.664 5.873 0.706 ;
      RECT 5.527 0.664 5.569 0.706 ;
      RECT 5.679 0.664 5.721 0.706 ;
      RECT 4.767 0.664 4.809 0.706 ;
      RECT 5.223 0.664 5.265 0.706 ;
      RECT 4.919 0.664 4.961 0.706 ;
      RECT 0.587 0.151 0.629 0.193 ;
      RECT 0.587 1.027 0.629 1.069 ;
      RECT 0.587 0.427 0.629 0.469 ;
      RECT 0.587 0.335 0.629 0.377 ;
      RECT 0.587 1.119 0.629 1.161 ;
      RECT 0.587 1.027 0.629 1.069 ;
      RECT 0.587 0.335 0.629 0.377 ;
      RECT 0.587 1.487 0.629 1.529 ;
      RECT 0.587 0.243 0.629 0.285 ;
      RECT 0.891 1.027 0.933 1.069 ;
      RECT 0.587 1.487 0.629 1.529 ;
      RECT 0.587 1.395 0.629 1.437 ;
      RECT 0.587 0.151 0.629 0.193 ;
      RECT 0.587 1.119 0.629 1.161 ;
      RECT 0.587 1.395 0.629 1.437 ;
      RECT 0.587 1.211 0.629 1.253 ;
      RECT 0.891 1.487 0.933 1.529 ;
      RECT 0.587 1.211 0.629 1.253 ;
      RECT 0.587 1.303 0.629 1.345 ;
      RECT 0.587 1.303 0.629 1.345 ;
      RECT 0.891 1.303 0.933 1.345 ;
      RECT 0.891 1.303 0.933 1.345 ;
      RECT 0.891 1.487 0.933 1.529 ;
      RECT 0.891 1.211 0.933 1.253 ;
      RECT 0.891 1.211 0.933 1.253 ;
      RECT 0.891 1.395 0.933 1.437 ;
      RECT 0.891 1.119 0.933 1.161 ;
      RECT 0.891 1.119 0.933 1.161 ;
      RECT 0.891 1.395 0.933 1.437 ;
      RECT 0.891 1.027 0.933 1.069 ;
      RECT 0.283 1.027 0.325 1.069 ;
      RECT 0.283 1.119 0.325 1.161 ;
      RECT 0.283 1.027 0.325 1.069 ;
      RECT 0.283 1.487 0.325 1.529 ;
      RECT 0.283 1.487 0.325 1.529 ;
      RECT 0.283 1.395 0.325 1.437 ;
      RECT 0.283 1.119 0.325 1.161 ;
      RECT 0.283 1.395 0.325 1.437 ;
      RECT 0.283 1.211 0.325 1.253 ;
      RECT 0.283 1.211 0.325 1.253 ;
      RECT 0.283 1.303 0.325 1.345 ;
      RECT 0.283 1.303 0.325 1.345 ;
      RECT 0.283 0.151 0.325 0.193 ;
      RECT 0.283 0.427 0.325 0.469 ;
      RECT 0.283 0.335 0.325 0.377 ;
      RECT 0.283 0.335 0.325 0.377 ;
      RECT 0.283 0.243 0.325 0.285 ;
      RECT 0.283 0.151 0.325 0.193 ;
      RECT 0.891 0.151 0.933 0.193 ;
      RECT 0.891 0.427 0.933 0.469 ;
      RECT 0.891 0.335 0.933 0.377 ;
      RECT 0.891 0.335 0.933 0.377 ;
      RECT 0.891 0.243 0.933 0.285 ;
      RECT 0.891 0.151 0.933 0.193 ;
      RECT 3.551 0.664 3.593 0.706 ;
      RECT 3.247 0.664 3.289 0.706 ;
      RECT 3.399 0.664 3.441 0.706 ;
      RECT 2.487 0.664 2.529 0.706 ;
      RECT 2.943 0.664 2.985 0.706 ;
      RECT 2.639 0.664 2.681 0.706 ;
      RECT 2.791 0.664 2.833 0.706 ;
      RECT 5.071 0.664 5.113 0.706 ;
      RECT 3.095 0.664 3.137 0.706 ;
      RECT 2.031 0.664 2.073 0.706 ;
      RECT 2.183 0.664 2.225 0.706 ;
      RECT 1.879 0.664 1.921 0.706 ;
      RECT 1.727 0.664 1.769 0.706 ;
      RECT 1.575 0.664 1.617 0.706 ;
      RECT 2.335 0.664 2.377 0.706 ;
      RECT 1.271 0.664 1.313 0.706 ;
      RECT 1.423 0.664 1.465 0.706 ;
    LAYER PO ;
      RECT 0.061 0.069 0.091 1.606 ;
      RECT 0.517 0.069 0.547 1.606 ;
      RECT 0.669 0.069 0.699 1.606 ;
      RECT 0.821 0.069 0.851 1.606 ;
      RECT 0.365 0.069 0.395 1.606 ;
      RECT 0.213 0.069 0.243 1.606 ;
      RECT 0.973 0.069 1.003 1.606 ;
      RECT 6.293 0.069 6.323 1.606 ;
      RECT 6.141 0.069 6.171 1.606 ;
      RECT 5.989 0.069 6.019 1.606 ;
      RECT 5.837 0.069 5.867 1.606 ;
      RECT 5.533 0.069 5.563 1.606 ;
      RECT 5.685 0.069 5.715 1.606 ;
      RECT 5.229 0.069 5.259 1.606 ;
      RECT 5.381 0.069 5.411 1.606 ;
      RECT 5.077 0.069 5.107 1.606 ;
      RECT 4.925 0.069 4.955 1.606 ;
      RECT 4.773 0.069 4.803 1.606 ;
      RECT 4.621 0.069 4.651 1.606 ;
      RECT 4.317 0.069 4.347 1.606 ;
      RECT 4.469 0.069 4.499 1.606 ;
      RECT 3.709 0.069 3.739 1.606 ;
      RECT 3.861 0.069 3.891 1.606 ;
      RECT 3.557 0.069 3.587 1.606 ;
      RECT 4.013 0.069 4.043 1.606 ;
      RECT 4.165 0.069 4.195 1.606 ;
      RECT 2.341 0.069 2.371 1.606 ;
      RECT 2.493 0.069 2.523 1.606 ;
      RECT 2.645 0.069 2.675 1.606 ;
      RECT 3.253 0.069 3.283 1.606 ;
      RECT 3.101 0.069 3.131 1.606 ;
      RECT 2.949 0.069 2.979 1.606 ;
      RECT 2.797 0.069 2.827 1.606 ;
      RECT 3.405 0.069 3.435 1.606 ;
      RECT 2.189 0.069 2.219 1.606 ;
      RECT 2.037 0.069 2.067 1.606 ;
      RECT 1.885 0.069 1.915 1.606 ;
      RECT 1.125 0.069 1.155 1.606 ;
      RECT 1.277 0.069 1.307 1.606 ;
      RECT 1.733 0.069 1.763 1.606 ;
      RECT 1.581 0.069 1.611 1.606 ;
      RECT 1.429 0.069 1.459 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 6.499 1.773 ;
  END
END NBUFFX32_RVT

MACRO IBUFFX16_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.952 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.664 0.401 0.706 ;
      LAYER M1 ;
        RECT 0.249 0.71 0.362 0.815 ;
        RECT 0.249 0.66 0.436 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.195 0.151 1.237 0.193 ;
        RECT 1.499 0.151 1.541 0.193 ;
        RECT 1.803 0.151 1.845 0.193 ;
        RECT 2.107 0.151 2.149 0.193 ;
        RECT 2.715 0.151 2.757 0.193 ;
        RECT 3.019 0.151 3.061 0.193 ;
        RECT 3.323 0.151 3.365 0.193 ;
        RECT 3.627 0.151 3.669 0.193 ;
        RECT 2.411 0.152 2.453 0.194 ;
        RECT 1.195 0.243 1.237 0.285 ;
        RECT 1.499 0.243 1.541 0.285 ;
        RECT 1.803 0.243 1.845 0.285 ;
        RECT 2.107 0.243 2.149 0.285 ;
        RECT 2.715 0.243 2.757 0.285 ;
        RECT 3.019 0.243 3.061 0.285 ;
        RECT 3.323 0.243 3.365 0.285 ;
        RECT 3.627 0.243 3.669 0.285 ;
        RECT 2.411 0.244 2.453 0.286 ;
        RECT 1.195 0.335 1.237 0.377 ;
        RECT 1.499 0.335 1.541 0.377 ;
        RECT 1.803 0.335 1.845 0.377 ;
        RECT 2.107 0.335 2.149 0.377 ;
        RECT 2.715 0.335 2.757 0.377 ;
        RECT 3.019 0.335 3.061 0.377 ;
        RECT 3.323 0.335 3.365 0.377 ;
        RECT 3.627 0.335 3.669 0.377 ;
        RECT 2.411 0.336 2.453 0.378 ;
        RECT 1.195 0.427 1.237 0.469 ;
        RECT 1.499 0.427 1.541 0.469 ;
        RECT 1.803 0.427 1.845 0.469 ;
        RECT 2.107 0.427 2.149 0.469 ;
        RECT 2.715 0.427 2.757 0.469 ;
        RECT 3.019 0.427 3.061 0.469 ;
        RECT 3.323 0.427 3.365 0.469 ;
        RECT 3.627 0.427 3.669 0.469 ;
        RECT 2.411 0.428 2.453 0.47 ;
        RECT 1.195 1.027 1.237 1.069 ;
        RECT 1.499 1.027 1.541 1.069 ;
        RECT 1.803 1.027 1.845 1.069 ;
        RECT 2.107 1.027 2.149 1.069 ;
        RECT 2.715 1.027 2.757 1.069 ;
        RECT 3.019 1.027 3.061 1.069 ;
        RECT 3.323 1.027 3.365 1.069 ;
        RECT 3.627 1.027 3.669 1.069 ;
        RECT 2.411 1.028 2.453 1.07 ;
        RECT 1.195 1.119 1.237 1.161 ;
        RECT 1.499 1.119 1.541 1.161 ;
        RECT 1.803 1.119 1.845 1.161 ;
        RECT 2.107 1.119 2.149 1.161 ;
        RECT 2.715 1.119 2.757 1.161 ;
        RECT 3.019 1.119 3.061 1.161 ;
        RECT 3.323 1.119 3.365 1.161 ;
        RECT 3.627 1.119 3.669 1.161 ;
        RECT 2.411 1.12 2.453 1.162 ;
        RECT 1.195 1.211 1.237 1.253 ;
        RECT 1.499 1.211 1.541 1.253 ;
        RECT 1.803 1.211 1.845 1.253 ;
        RECT 2.107 1.211 2.149 1.253 ;
        RECT 2.715 1.211 2.757 1.253 ;
        RECT 3.019 1.211 3.061 1.253 ;
        RECT 3.323 1.211 3.365 1.253 ;
        RECT 3.627 1.211 3.669 1.253 ;
        RECT 2.411 1.212 2.453 1.254 ;
        RECT 1.195 1.303 1.237 1.345 ;
        RECT 1.499 1.303 1.541 1.345 ;
        RECT 1.803 1.303 1.845 1.345 ;
        RECT 2.107 1.303 2.149 1.345 ;
        RECT 2.715 1.303 2.757 1.345 ;
        RECT 3.019 1.303 3.061 1.345 ;
        RECT 3.323 1.303 3.365 1.345 ;
        RECT 3.627 1.303 3.669 1.345 ;
        RECT 2.411 1.304 2.453 1.346 ;
        RECT 1.195 1.395 1.237 1.437 ;
        RECT 1.499 1.395 1.541 1.437 ;
        RECT 1.803 1.395 1.845 1.437 ;
        RECT 2.107 1.395 2.149 1.437 ;
        RECT 2.715 1.395 2.757 1.437 ;
        RECT 3.019 1.395 3.061 1.437 ;
        RECT 3.323 1.395 3.365 1.437 ;
        RECT 3.627 1.395 3.669 1.437 ;
        RECT 2.411 1.396 2.453 1.438 ;
        RECT 1.195 1.487 1.237 1.529 ;
        RECT 1.499 1.487 1.541 1.529 ;
        RECT 1.803 1.487 1.845 1.529 ;
        RECT 2.107 1.487 2.149 1.529 ;
        RECT 2.715 1.487 2.757 1.529 ;
        RECT 3.019 1.487 3.061 1.529 ;
        RECT 3.323 1.487 3.365 1.529 ;
        RECT 3.627 1.487 3.669 1.529 ;
        RECT 2.411 1.488 2.453 1.53 ;
      LAYER M1 ;
        RECT 2.407 0.942 2.457 1.565 ;
        RECT 1.191 0.942 1.241 1.564 ;
        RECT 1.495 0.942 1.545 1.564 ;
        RECT 1.799 0.942 1.849 1.564 ;
        RECT 2.103 0.942 2.153 1.564 ;
        RECT 2.711 0.942 2.761 1.564 ;
        RECT 3.015 0.942 3.065 1.564 ;
        RECT 3.319 0.942 3.369 1.564 ;
        RECT 3.623 0.942 3.673 1.564 ;
        RECT 1.191 0.892 3.732 0.942 ;
        RECT 3.682 0.663 3.732 0.892 ;
        RECT 3.682 0.587 3.855 0.663 ;
        RECT 1.191 0.537 3.855 0.587 ;
        RECT 1.191 0.116 1.241 0.537 ;
        RECT 1.495 0.116 1.545 0.537 ;
        RECT 1.799 0.116 1.849 0.537 ;
        RECT 2.103 0.116 2.153 0.537 ;
        RECT 2.407 0.117 2.457 0.537 ;
        RECT 2.711 0.116 2.761 0.537 ;
        RECT 3.015 0.116 3.065 0.537 ;
        RECT 3.319 0.116 3.369 0.537 ;
        RECT 3.623 0.116 3.673 0.537 ;
    END
    ANTENNADIFFAREA 1.2904 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.435 1.027 0.477 1.069 ;
        RECT 0.739 1.027 0.781 1.069 ;
        RECT 1.043 1.027 1.085 1.069 ;
        RECT 1.347 1.027 1.389 1.069 ;
        RECT 1.651 1.027 1.693 1.069 ;
        RECT 1.955 1.027 1.997 1.069 ;
        RECT 2.259 1.027 2.301 1.069 ;
        RECT 2.563 1.027 2.605 1.069 ;
        RECT 2.867 1.027 2.909 1.069 ;
        RECT 3.171 1.027 3.213 1.069 ;
        RECT 3.475 1.027 3.517 1.069 ;
        RECT 0.435 1.119 0.477 1.161 ;
        RECT 0.739 1.119 0.781 1.161 ;
        RECT 1.043 1.119 1.085 1.161 ;
        RECT 1.347 1.119 1.389 1.161 ;
        RECT 1.651 1.119 1.693 1.161 ;
        RECT 1.955 1.119 1.997 1.161 ;
        RECT 2.259 1.119 2.301 1.161 ;
        RECT 2.563 1.119 2.605 1.161 ;
        RECT 2.867 1.119 2.909 1.161 ;
        RECT 3.171 1.119 3.213 1.161 ;
        RECT 3.475 1.119 3.517 1.161 ;
        RECT 0.435 1.211 0.477 1.253 ;
        RECT 0.739 1.211 0.781 1.253 ;
        RECT 1.043 1.211 1.085 1.253 ;
        RECT 1.347 1.211 1.389 1.253 ;
        RECT 1.651 1.211 1.693 1.253 ;
        RECT 1.955 1.211 1.997 1.253 ;
        RECT 2.259 1.211 2.301 1.253 ;
        RECT 2.563 1.211 2.605 1.253 ;
        RECT 2.867 1.211 2.909 1.253 ;
        RECT 3.171 1.211 3.213 1.253 ;
        RECT 3.475 1.211 3.517 1.253 ;
        RECT 0.435 1.303 0.477 1.345 ;
        RECT 0.739 1.303 0.781 1.345 ;
        RECT 1.043 1.303 1.085 1.345 ;
        RECT 1.347 1.303 1.389 1.345 ;
        RECT 1.651 1.303 1.693 1.345 ;
        RECT 1.955 1.303 1.997 1.345 ;
        RECT 2.259 1.303 2.301 1.345 ;
        RECT 2.563 1.303 2.605 1.345 ;
        RECT 2.867 1.303 2.909 1.345 ;
        RECT 3.171 1.303 3.213 1.345 ;
        RECT 3.475 1.303 3.517 1.345 ;
        RECT 0.435 1.395 0.477 1.437 ;
        RECT 0.739 1.395 0.781 1.437 ;
        RECT 1.043 1.395 1.085 1.437 ;
        RECT 1.347 1.395 1.389 1.437 ;
        RECT 1.651 1.395 1.693 1.437 ;
        RECT 1.955 1.395 1.997 1.437 ;
        RECT 2.259 1.395 2.301 1.437 ;
        RECT 2.563 1.395 2.605 1.437 ;
        RECT 2.867 1.395 2.909 1.437 ;
        RECT 3.171 1.395 3.213 1.437 ;
        RECT 3.475 1.395 3.517 1.437 ;
        RECT 0.435 1.487 0.477 1.529 ;
        RECT 0.739 1.487 0.781 1.529 ;
        RECT 1.043 1.487 1.085 1.529 ;
        RECT 1.347 1.487 1.389 1.529 ;
        RECT 1.651 1.487 1.693 1.529 ;
        RECT 1.955 1.487 1.997 1.529 ;
        RECT 2.259 1.487 2.301 1.529 ;
        RECT 2.563 1.487 2.605 1.529 ;
        RECT 2.867 1.487 2.909 1.529 ;
        RECT 3.171 1.487 3.213 1.529 ;
        RECT 3.475 1.487 3.517 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
        RECT 3.095 1.651 3.137 1.693 ;
        RECT 3.247 1.651 3.289 1.693 ;
        RECT 3.399 1.651 3.441 1.693 ;
        RECT 3.551 1.651 3.593 1.693 ;
        RECT 3.703 1.651 3.745 1.693 ;
        RECT 3.855 1.651 3.897 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 3.952 1.702 ;
        RECT 0.431 0.992 0.481 1.642 ;
        RECT 0.735 0.992 0.785 1.642 ;
        RECT 1.039 0.992 1.089 1.642 ;
        RECT 1.343 0.992 1.393 1.642 ;
        RECT 1.647 0.992 1.697 1.642 ;
        RECT 1.951 0.992 2.001 1.642 ;
        RECT 2.255 0.992 2.305 1.642 ;
        RECT 2.559 0.992 2.609 1.642 ;
        RECT 2.863 0.992 2.913 1.642 ;
        RECT 3.167 0.992 3.217 1.642 ;
        RECT 3.471 0.992 3.521 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 3.399 -0.021 3.441 0.021 ;
        RECT 3.551 -0.021 3.593 0.021 ;
        RECT 3.703 -0.021 3.745 0.021 ;
        RECT 3.855 -0.021 3.897 0.021 ;
        RECT 0.435 0.149 0.477 0.191 ;
        RECT 0.739 0.149 0.781 0.191 ;
        RECT 1.043 0.149 1.085 0.191 ;
        RECT 1.347 0.149 1.389 0.191 ;
        RECT 1.651 0.149 1.693 0.191 ;
        RECT 1.955 0.149 1.997 0.191 ;
        RECT 2.259 0.149 2.301 0.191 ;
        RECT 2.563 0.149 2.605 0.191 ;
        RECT 2.867 0.149 2.909 0.191 ;
        RECT 3.171 0.149 3.213 0.191 ;
        RECT 3.475 0.149 3.517 0.191 ;
        RECT 0.435 0.241 0.477 0.283 ;
        RECT 0.739 0.241 0.781 0.283 ;
        RECT 1.043 0.241 1.085 0.283 ;
        RECT 1.347 0.241 1.389 0.283 ;
        RECT 1.651 0.241 1.693 0.283 ;
        RECT 1.955 0.241 1.997 0.283 ;
        RECT 2.259 0.241 2.301 0.283 ;
        RECT 2.563 0.241 2.605 0.283 ;
        RECT 2.867 0.241 2.909 0.283 ;
        RECT 3.171 0.241 3.213 0.283 ;
        RECT 3.475 0.241 3.517 0.283 ;
        RECT 0.435 0.333 0.477 0.375 ;
        RECT 0.739 0.333 0.781 0.375 ;
        RECT 1.043 0.333 1.085 0.375 ;
        RECT 1.347 0.333 1.389 0.375 ;
        RECT 1.651 0.333 1.693 0.375 ;
        RECT 1.955 0.333 1.997 0.375 ;
        RECT 2.259 0.333 2.301 0.375 ;
        RECT 2.563 0.333 2.605 0.375 ;
        RECT 2.867 0.333 2.909 0.375 ;
        RECT 3.171 0.333 3.213 0.375 ;
        RECT 3.475 0.333 3.517 0.375 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.41 ;
        RECT 0.735 0.03 0.785 0.41 ;
        RECT 1.039 0.03 1.089 0.41 ;
        RECT 1.343 0.03 1.393 0.41 ;
        RECT 1.647 0.03 1.697 0.41 ;
        RECT 1.951 0.03 2.001 0.41 ;
        RECT 2.255 0.03 2.305 0.41 ;
        RECT 2.559 0.03 2.609 0.41 ;
        RECT 2.863 0.03 2.913 0.41 ;
        RECT 3.167 0.03 3.217 0.41 ;
        RECT 3.471 0.03 3.521 0.41 ;
        RECT 0 -0.03 3.952 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.891 1.119 0.933 1.161 ;
      RECT 0.891 1.395 0.933 1.437 ;
      RECT 0.891 1.211 0.933 1.253 ;
      RECT 0.283 1.487 0.325 1.529 ;
      RECT 0.283 1.487 0.325 1.529 ;
      RECT 2.943 0.664 2.985 0.706 ;
      RECT 2.639 0.664 2.681 0.706 ;
      RECT 2.791 0.664 2.833 0.706 ;
      RECT 0.283 1.211 0.325 1.253 ;
      RECT 0.283 0.427 0.325 0.469 ;
      RECT 0.891 1.211 0.933 1.253 ;
      RECT 0.815 0.664 0.857 0.706 ;
      RECT 0.283 1.395 0.325 1.437 ;
      RECT 0.891 1.303 0.933 1.345 ;
      RECT 0.663 0.664 0.705 0.706 ;
      RECT 0.891 1.303 0.933 1.345 ;
      RECT 0.283 0.243 0.325 0.285 ;
      RECT 0.283 0.151 0.325 0.193 ;
      RECT 0.283 0.151 0.325 0.193 ;
      RECT 0.283 1.303 0.325 1.345 ;
      RECT 0.283 0.335 0.325 0.377 ;
      RECT 0.283 1.303 0.325 1.345 ;
      RECT 0.283 0.335 0.325 0.377 ;
      RECT 0.587 1.027 0.629 1.069 ;
      RECT 0.587 1.119 0.629 1.161 ;
      RECT 0.587 1.027 0.629 1.069 ;
      RECT 0.587 1.487 0.629 1.529 ;
      RECT 0.587 1.487 0.629 1.529 ;
      RECT 0.587 1.395 0.629 1.437 ;
      RECT 0.587 1.119 0.629 1.161 ;
      RECT 0.587 1.395 0.629 1.437 ;
      RECT 0.587 1.211 0.629 1.253 ;
      RECT 0.587 1.211 0.629 1.253 ;
      RECT 0.587 1.303 0.629 1.345 ;
      RECT 0.587 1.303 0.629 1.345 ;
      RECT 0.587 0.151 0.629 0.193 ;
      RECT 0.587 0.427 0.629 0.469 ;
      RECT 0.587 0.335 0.629 0.377 ;
      RECT 0.587 0.335 0.629 0.377 ;
      RECT 0.587 0.243 0.629 0.285 ;
      RECT 0.587 0.151 0.629 0.193 ;
      RECT 3.095 0.664 3.137 0.706 ;
      RECT 3.551 0.664 3.593 0.706 ;
      RECT 3.247 0.664 3.289 0.706 ;
      RECT 3.399 0.664 3.441 0.706 ;
      RECT 0.283 1.119 0.325 1.161 ;
      RECT 0.891 0.151 0.933 0.193 ;
      RECT 0.891 1.027 0.933 1.069 ;
      RECT 0.283 1.395 0.325 1.437 ;
      RECT 0.891 0.427 0.933 0.469 ;
      RECT 0.891 0.335 0.933 0.377 ;
      RECT 0.891 1.119 0.933 1.161 ;
      RECT 0.283 1.027 0.325 1.069 ;
      RECT 0.283 1.119 0.325 1.161 ;
      RECT 0.891 1.027 0.933 1.069 ;
      RECT 0.283 1.027 0.325 1.069 ;
      RECT 0.891 0.335 0.933 0.377 ;
      RECT 0.891 1.487 0.933 1.529 ;
      RECT 0.891 0.243 0.933 0.285 ;
      RECT 0.891 1.487 0.933 1.529 ;
      RECT 0.283 1.211 0.325 1.253 ;
      RECT 0.891 1.395 0.933 1.437 ;
      RECT 0.891 0.151 0.933 0.193 ;
      RECT 2.335 0.664 2.377 0.706 ;
      RECT 2.487 0.664 2.529 0.706 ;
      RECT 1.271 0.664 1.313 0.706 ;
      RECT 0.967 0.664 1.009 0.706 ;
      RECT 1.423 0.664 1.465 0.706 ;
      RECT 2.031 0.664 2.073 0.706 ;
      RECT 2.183 0.664 2.225 0.706 ;
      RECT 1.879 0.664 1.921 0.706 ;
      RECT 1.727 0.664 1.769 0.706 ;
      RECT 1.575 0.664 1.617 0.706 ;
    LAYER M1 ;
      RECT 1.094 0.66 3.628 0.71 ;
      RECT 0.583 0.942 0.633 1.564 ;
      RECT 0.583 0.116 0.633 0.537 ;
      RECT 0.887 0.942 0.937 1.564 ;
      RECT 0.887 0.116 0.937 0.537 ;
      RECT 0.583 0.537 1.141 0.587 ;
      RECT 1.091 0.605 1.144 0.633 ;
      RECT 1.094 0.633 1.144 0.66 ;
      RECT 1.091 0.587 1.141 0.605 ;
      RECT 1.094 0.71 1.144 0.842 ;
      RECT 1.09 0.874 1.14 0.892 ;
      RECT 1.09 0.842 1.144 0.874 ;
      RECT 0.583 0.892 1.14 0.942 ;
      RECT 0.487 0.66 1.044 0.71 ;
      RECT 0.279 0.942 0.329 1.564 ;
      RECT 0.279 0.116 0.329 0.537 ;
      RECT 0.279 0.892 0.533 0.942 ;
      RECT 0.483 0.832 0.537 0.87 ;
      RECT 0.279 0.537 0.533 0.587 ;
      RECT 0.487 0.71 0.537 0.832 ;
      RECT 0.483 0.87 0.533 0.892 ;
      RECT 0.487 0.642 0.537 0.66 ;
      RECT 0.483 0.587 0.533 0.607 ;
      RECT 0.483 0.607 0.537 0.642 ;
    LAYER PO ;
      RECT 3.861 0.069 3.891 1.606 ;
      RECT 3.557 0.069 3.587 1.606 ;
      RECT 2.341 0.069 2.371 1.606 ;
      RECT 2.493 0.069 2.523 1.606 ;
      RECT 2.645 0.069 2.675 1.606 ;
      RECT 3.253 0.069 3.283 1.606 ;
      RECT 3.101 0.069 3.131 1.606 ;
      RECT 2.949 0.069 2.979 1.606 ;
      RECT 2.797 0.069 2.827 1.606 ;
      RECT 3.405 0.069 3.435 1.606 ;
      RECT 2.189 0.069 2.219 1.606 ;
      RECT 2.037 0.069 2.067 1.606 ;
      RECT 1.885 0.069 1.915 1.606 ;
      RECT 1.125 0.069 1.155 1.606 ;
      RECT 1.277 0.069 1.307 1.606 ;
      RECT 1.733 0.069 1.763 1.606 ;
      RECT 1.581 0.069 1.611 1.606 ;
      RECT 1.429 0.069 1.459 1.606 ;
      RECT 0.061 0.071 0.091 1.606 ;
      RECT 0.821 0.069 0.851 1.606 ;
      RECT 0.973 0.069 1.003 1.606 ;
      RECT 0.365 0.069 0.395 1.606 ;
      RECT 0.669 0.069 0.699 1.606 ;
      RECT 0.213 0.071 0.243 1.606 ;
      RECT 0.517 0.071 0.547 1.606 ;
      RECT 3.709 0.069 3.739 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 4.067 1.773 ;
  END
END IBUFFX16_RVT

MACRO IBUFFX2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.664 0.401 0.706 ;
      LAYER M1 ;
        RECT 0.249 0.71 0.362 0.815 ;
        RECT 0.249 0.66 0.436 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0186 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.891 0.151 0.933 0.193 ;
        RECT 1.195 0.151 1.237 0.193 ;
        RECT 0.891 0.243 0.933 0.285 ;
        RECT 1.195 0.243 1.237 0.285 ;
        RECT 0.891 0.335 0.933 0.377 ;
        RECT 1.195 0.335 1.237 0.377 ;
        RECT 0.891 0.427 0.933 0.469 ;
        RECT 1.195 0.427 1.237 0.469 ;
        RECT 0.891 1.027 0.933 1.069 ;
        RECT 1.195 1.027 1.237 1.069 ;
        RECT 0.891 1.119 0.933 1.161 ;
        RECT 1.195 1.119 1.237 1.161 ;
        RECT 0.891 1.211 0.933 1.253 ;
        RECT 1.195 1.211 1.237 1.253 ;
        RECT 0.891 1.303 0.933 1.345 ;
        RECT 1.195 1.303 1.237 1.345 ;
        RECT 0.891 1.395 0.933 1.437 ;
        RECT 1.195 1.395 1.237 1.437 ;
        RECT 0.891 1.487 0.933 1.529 ;
        RECT 1.195 1.487 1.237 1.529 ;
      LAYER M1 ;
        RECT 0.887 0.942 0.937 1.564 ;
        RECT 1.191 0.942 1.241 1.564 ;
        RECT 0.887 0.892 1.297 0.942 ;
        RECT 1.247 0.663 1.297 0.892 ;
        RECT 1.247 0.587 1.423 0.663 ;
        RECT 0.887 0.537 1.423 0.587 ;
        RECT 0.887 0.116 0.937 0.537 ;
        RECT 1.191 0.116 1.241 0.537 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 0.9 0.325 0.942 ;
        RECT 0.587 0.929 0.629 0.971 ;
        RECT 0.283 0.992 0.325 1.034 ;
        RECT 0.587 1.022 0.629 1.064 ;
        RECT 1.043 1.027 1.085 1.069 ;
        RECT 0.283 1.084 0.325 1.126 ;
        RECT 0.587 1.114 0.629 1.156 ;
        RECT 1.043 1.119 1.085 1.161 ;
        RECT 1.043 1.211 1.085 1.253 ;
        RECT 1.043 1.303 1.085 1.345 ;
        RECT 1.043 1.395 1.085 1.437 ;
        RECT 1.043 1.487 1.085 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.52 1.702 ;
        RECT 0.279 0.865 0.329 1.642 ;
        RECT 0.583 0.893 0.633 1.642 ;
        RECT 1.039 0.992 1.089 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.043 0.149 1.085 0.191 ;
        RECT 1.043 0.241 1.085 0.283 ;
        RECT 0.587 0.305 0.629 0.347 ;
        RECT 1.043 0.333 1.085 0.375 ;
        RECT 0.283 0.378 0.325 0.42 ;
        RECT 0.587 0.397 0.629 0.439 ;
        RECT 0.283 0.47 0.325 0.512 ;
        RECT 0.587 0.489 0.629 0.531 ;
      LAYER M1 ;
        RECT 0.279 0.03 0.329 0.56 ;
        RECT 0.583 0.03 0.633 0.554 ;
        RECT 1.039 0.03 1.089 0.41 ;
        RECT 0 -0.03 1.52 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.663 0.664 0.705 0.706 ;
      RECT 0.739 0.93 0.781 0.972 ;
      RECT 0.967 0.664 1.009 0.706 ;
      RECT 0.739 1.114 0.781 1.156 ;
      RECT 0.739 1.022 0.781 1.064 ;
      RECT 0.739 0.93 0.781 0.972 ;
      RECT 0.739 0.489 0.781 0.531 ;
      RECT 0.739 0.397 0.781 0.439 ;
      RECT 0.739 0.397 0.781 0.439 ;
      RECT 1.119 0.664 1.161 0.706 ;
      RECT 0.739 1.022 0.781 1.064 ;
      RECT 0.739 1.114 0.781 1.156 ;
      RECT 0.435 1.086 0.477 1.128 ;
      RECT 0.435 0.81 0.477 0.852 ;
      RECT 0.435 0.902 0.477 0.944 ;
      RECT 0.435 0.994 0.477 1.036 ;
      RECT 0.435 1.086 0.477 1.128 ;
      RECT 0.435 0.81 0.477 0.852 ;
      RECT 0.435 0.483 0.477 0.525 ;
      RECT 0.435 0.994 0.477 1.036 ;
      RECT 0.435 0.391 0.477 0.433 ;
      RECT 0.435 0.902 0.477 0.944 ;
      RECT 0.739 0.835 0.781 0.877 ;
      RECT 0.435 0.391 0.477 0.433 ;
      RECT 0.739 0.305 0.781 0.347 ;
      RECT 0.739 0.835 0.781 0.877 ;
    LAYER M1 ;
      RECT 0.487 0.66 0.74 0.71 ;
      RECT 0.431 0.362 0.481 0.532 ;
      RECT 0.431 0.532 0.533 0.582 ;
      RECT 0.487 0.71 0.537 0.775 ;
      RECT 0.431 0.775 0.537 0.825 ;
      RECT 0.431 0.825 0.481 1.165 ;
      RECT 0.487 0.63 0.537 0.66 ;
      RECT 0.483 0.582 0.533 0.607 ;
      RECT 0.483 0.607 0.537 0.63 ;
      RECT 0.791 0.66 1.196 0.71 ;
      RECT 0.735 0.776 0.841 0.826 ;
      RECT 0.735 0.826 0.785 1.191 ;
      RECT 0.735 0.532 0.837 0.582 ;
      RECT 0.791 0.71 0.841 0.776 ;
      RECT 0.735 0.285 0.785 0.532 ;
      RECT 0.791 0.641 0.841 0.66 ;
      RECT 0.787 0.582 0.837 0.607 ;
      RECT 0.787 0.607 0.841 0.641 ;
    LAYER PO ;
      RECT 0.061 0.069 0.091 1.606 ;
      RECT 0.213 0.069 0.243 1.606 ;
      RECT 0.365 0.071 0.395 1.606 ;
      RECT 0.669 0.069 0.699 1.606 ;
      RECT 0.517 0.071 0.547 1.606 ;
      RECT 0.821 0.071 0.851 1.606 ;
      RECT 0.973 0.069 1.003 1.606 ;
      RECT 1.429 0.071 1.459 1.606 ;
      RECT 1.277 0.071 1.307 1.606 ;
      RECT 1.125 0.069 1.155 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.635 1.773 ;
  END
END IBUFFX2_RVT

MACRO IBUFFX32_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 6.992 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.664 0.401 0.706 ;
        RECT 0.511 0.664 0.553 0.706 ;
      LAYER M1 ;
        RECT 0.249 0.71 0.362 0.815 ;
        RECT 0.249 0.66 0.588 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0732 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.803 0.151 1.845 0.193 ;
        RECT 2.107 0.151 2.149 0.193 ;
        RECT 2.411 0.151 2.453 0.193 ;
        RECT 2.715 0.151 2.757 0.193 ;
        RECT 3.323 0.151 3.365 0.193 ;
        RECT 3.627 0.151 3.669 0.193 ;
        RECT 3.931 0.151 3.973 0.193 ;
        RECT 4.235 0.151 4.277 0.193 ;
        RECT 4.539 0.151 4.581 0.193 ;
        RECT 4.843 0.151 4.885 0.193 ;
        RECT 5.147 0.151 5.189 0.193 ;
        RECT 5.451 0.151 5.493 0.193 ;
        RECT 5.755 0.151 5.797 0.193 ;
        RECT 6.059 0.151 6.101 0.193 ;
        RECT 6.363 0.151 6.405 0.193 ;
        RECT 6.667 0.151 6.709 0.193 ;
        RECT 3.019 0.152 3.061 0.194 ;
        RECT 1.803 0.243 1.845 0.285 ;
        RECT 2.107 0.243 2.149 0.285 ;
        RECT 2.411 0.243 2.453 0.285 ;
        RECT 2.715 0.243 2.757 0.285 ;
        RECT 3.323 0.243 3.365 0.285 ;
        RECT 3.627 0.243 3.669 0.285 ;
        RECT 3.931 0.243 3.973 0.285 ;
        RECT 4.235 0.243 4.277 0.285 ;
        RECT 4.539 0.243 4.581 0.285 ;
        RECT 4.843 0.243 4.885 0.285 ;
        RECT 5.147 0.243 5.189 0.285 ;
        RECT 5.451 0.243 5.493 0.285 ;
        RECT 5.755 0.243 5.797 0.285 ;
        RECT 6.059 0.243 6.101 0.285 ;
        RECT 6.363 0.243 6.405 0.285 ;
        RECT 6.667 0.243 6.709 0.285 ;
        RECT 3.019 0.244 3.061 0.286 ;
        RECT 1.803 0.335 1.845 0.377 ;
        RECT 2.107 0.335 2.149 0.377 ;
        RECT 2.411 0.335 2.453 0.377 ;
        RECT 2.715 0.335 2.757 0.377 ;
        RECT 3.323 0.335 3.365 0.377 ;
        RECT 3.627 0.335 3.669 0.377 ;
        RECT 3.931 0.335 3.973 0.377 ;
        RECT 4.235 0.335 4.277 0.377 ;
        RECT 4.539 0.335 4.581 0.377 ;
        RECT 4.843 0.335 4.885 0.377 ;
        RECT 5.147 0.335 5.189 0.377 ;
        RECT 5.451 0.335 5.493 0.377 ;
        RECT 5.755 0.335 5.797 0.377 ;
        RECT 6.059 0.335 6.101 0.377 ;
        RECT 6.363 0.335 6.405 0.377 ;
        RECT 6.667 0.335 6.709 0.377 ;
        RECT 3.019 0.336 3.061 0.378 ;
        RECT 1.803 0.427 1.845 0.469 ;
        RECT 2.107 0.427 2.149 0.469 ;
        RECT 2.411 0.427 2.453 0.469 ;
        RECT 2.715 0.427 2.757 0.469 ;
        RECT 3.323 0.427 3.365 0.469 ;
        RECT 3.627 0.427 3.669 0.469 ;
        RECT 3.931 0.427 3.973 0.469 ;
        RECT 4.235 0.427 4.277 0.469 ;
        RECT 4.539 0.427 4.581 0.469 ;
        RECT 4.843 0.427 4.885 0.469 ;
        RECT 5.147 0.427 5.189 0.469 ;
        RECT 5.451 0.427 5.493 0.469 ;
        RECT 5.755 0.427 5.797 0.469 ;
        RECT 6.059 0.427 6.101 0.469 ;
        RECT 6.363 0.427 6.405 0.469 ;
        RECT 6.667 0.427 6.709 0.469 ;
        RECT 3.019 0.428 3.061 0.47 ;
        RECT 1.803 1.027 1.845 1.069 ;
        RECT 2.107 1.027 2.149 1.069 ;
        RECT 2.411 1.027 2.453 1.069 ;
        RECT 2.715 1.027 2.757 1.069 ;
        RECT 3.323 1.027 3.365 1.069 ;
        RECT 3.627 1.027 3.669 1.069 ;
        RECT 3.931 1.027 3.973 1.069 ;
        RECT 4.235 1.027 4.277 1.069 ;
        RECT 4.539 1.027 4.581 1.069 ;
        RECT 4.843 1.027 4.885 1.069 ;
        RECT 5.147 1.027 5.189 1.069 ;
        RECT 5.451 1.027 5.493 1.069 ;
        RECT 5.755 1.027 5.797 1.069 ;
        RECT 6.059 1.027 6.101 1.069 ;
        RECT 6.363 1.027 6.405 1.069 ;
        RECT 6.667 1.027 6.709 1.069 ;
        RECT 3.019 1.028 3.061 1.07 ;
        RECT 1.803 1.119 1.845 1.161 ;
        RECT 2.107 1.119 2.149 1.161 ;
        RECT 2.411 1.119 2.453 1.161 ;
        RECT 2.715 1.119 2.757 1.161 ;
        RECT 3.323 1.119 3.365 1.161 ;
        RECT 3.627 1.119 3.669 1.161 ;
        RECT 3.931 1.119 3.973 1.161 ;
        RECT 4.235 1.119 4.277 1.161 ;
        RECT 4.539 1.119 4.581 1.161 ;
        RECT 4.843 1.119 4.885 1.161 ;
        RECT 5.147 1.119 5.189 1.161 ;
        RECT 5.451 1.119 5.493 1.161 ;
        RECT 5.755 1.119 5.797 1.161 ;
        RECT 6.059 1.119 6.101 1.161 ;
        RECT 6.363 1.119 6.405 1.161 ;
        RECT 6.667 1.119 6.709 1.161 ;
        RECT 3.019 1.12 3.061 1.162 ;
        RECT 1.803 1.211 1.845 1.253 ;
        RECT 2.107 1.211 2.149 1.253 ;
        RECT 2.411 1.211 2.453 1.253 ;
        RECT 2.715 1.211 2.757 1.253 ;
        RECT 3.323 1.211 3.365 1.253 ;
        RECT 3.627 1.211 3.669 1.253 ;
        RECT 3.931 1.211 3.973 1.253 ;
        RECT 4.235 1.211 4.277 1.253 ;
        RECT 4.539 1.211 4.581 1.253 ;
        RECT 4.843 1.211 4.885 1.253 ;
        RECT 5.147 1.211 5.189 1.253 ;
        RECT 5.451 1.211 5.493 1.253 ;
        RECT 5.755 1.211 5.797 1.253 ;
        RECT 6.059 1.211 6.101 1.253 ;
        RECT 6.363 1.211 6.405 1.253 ;
        RECT 6.667 1.211 6.709 1.253 ;
        RECT 3.019 1.212 3.061 1.254 ;
        RECT 1.803 1.303 1.845 1.345 ;
        RECT 2.107 1.303 2.149 1.345 ;
        RECT 2.411 1.303 2.453 1.345 ;
        RECT 2.715 1.303 2.757 1.345 ;
        RECT 3.323 1.303 3.365 1.345 ;
        RECT 3.627 1.303 3.669 1.345 ;
        RECT 3.931 1.303 3.973 1.345 ;
        RECT 4.235 1.303 4.277 1.345 ;
        RECT 4.539 1.303 4.581 1.345 ;
        RECT 4.843 1.303 4.885 1.345 ;
        RECT 5.147 1.303 5.189 1.345 ;
        RECT 5.451 1.303 5.493 1.345 ;
        RECT 5.755 1.303 5.797 1.345 ;
        RECT 6.059 1.303 6.101 1.345 ;
        RECT 6.363 1.303 6.405 1.345 ;
        RECT 6.667 1.303 6.709 1.345 ;
        RECT 3.019 1.304 3.061 1.346 ;
        RECT 1.803 1.395 1.845 1.437 ;
        RECT 2.107 1.395 2.149 1.437 ;
        RECT 2.411 1.395 2.453 1.437 ;
        RECT 2.715 1.395 2.757 1.437 ;
        RECT 3.323 1.395 3.365 1.437 ;
        RECT 3.627 1.395 3.669 1.437 ;
        RECT 3.931 1.395 3.973 1.437 ;
        RECT 4.235 1.395 4.277 1.437 ;
        RECT 4.539 1.395 4.581 1.437 ;
        RECT 4.843 1.395 4.885 1.437 ;
        RECT 5.147 1.395 5.189 1.437 ;
        RECT 5.451 1.395 5.493 1.437 ;
        RECT 5.755 1.395 5.797 1.437 ;
        RECT 6.059 1.395 6.101 1.437 ;
        RECT 6.363 1.395 6.405 1.437 ;
        RECT 6.667 1.395 6.709 1.437 ;
        RECT 3.019 1.396 3.061 1.438 ;
        RECT 1.803 1.487 1.845 1.529 ;
        RECT 2.107 1.487 2.149 1.529 ;
        RECT 2.411 1.487 2.453 1.529 ;
        RECT 2.715 1.487 2.757 1.529 ;
        RECT 3.323 1.487 3.365 1.529 ;
        RECT 3.627 1.487 3.669 1.529 ;
        RECT 3.931 1.487 3.973 1.529 ;
        RECT 4.235 1.487 4.277 1.529 ;
        RECT 4.539 1.487 4.581 1.529 ;
        RECT 4.843 1.487 4.885 1.529 ;
        RECT 5.147 1.487 5.189 1.529 ;
        RECT 5.451 1.487 5.493 1.529 ;
        RECT 5.755 1.487 5.797 1.529 ;
        RECT 6.059 1.487 6.101 1.529 ;
        RECT 6.363 1.487 6.405 1.529 ;
        RECT 6.667 1.487 6.709 1.529 ;
        RECT 3.019 1.488 3.061 1.53 ;
      LAYER M1 ;
        RECT 4.535 0.942 4.585 1.564 ;
        RECT 4.839 0.942 4.889 1.564 ;
        RECT 5.143 0.942 5.193 1.564 ;
        RECT 5.447 0.942 5.497 1.564 ;
        RECT 5.751 0.942 5.801 1.564 ;
        RECT 6.055 0.942 6.105 1.564 ;
        RECT 6.359 0.942 6.409 1.564 ;
        RECT 6.663 0.942 6.713 1.564 ;
        RECT 6.722 0.663 6.772 0.892 ;
        RECT 1.799 0.892 6.772 0.942 ;
        RECT 3.015 0.942 3.065 1.565 ;
        RECT 1.799 0.942 1.849 1.564 ;
        RECT 2.103 0.942 2.153 1.564 ;
        RECT 2.407 0.942 2.457 1.564 ;
        RECT 2.711 0.942 2.761 1.564 ;
        RECT 3.319 0.942 3.369 1.564 ;
        RECT 3.623 0.942 3.673 1.564 ;
        RECT 3.927 0.942 3.977 1.564 ;
        RECT 4.231 0.942 4.281 1.564 ;
        RECT 6.722 0.587 6.895 0.663 ;
        RECT 1.799 0.537 6.895 0.587 ;
        RECT 4.535 0.116 4.585 0.537 ;
        RECT 4.839 0.116 4.889 0.537 ;
        RECT 5.143 0.116 5.193 0.537 ;
        RECT 5.447 0.116 5.497 0.537 ;
        RECT 5.751 0.116 5.801 0.537 ;
        RECT 6.055 0.116 6.105 0.537 ;
        RECT 6.359 0.116 6.409 0.537 ;
        RECT 6.663 0.116 6.713 0.537 ;
        RECT 1.799 0.116 1.849 0.537 ;
        RECT 2.103 0.116 2.153 0.537 ;
        RECT 2.407 0.116 2.457 0.537 ;
        RECT 2.711 0.116 2.761 0.537 ;
        RECT 3.015 0.117 3.065 0.537 ;
        RECT 3.319 0.116 3.369 0.537 ;
        RECT 3.623 0.116 3.673 0.537 ;
        RECT 3.927 0.116 3.977 0.537 ;
        RECT 4.231 0.116 4.281 0.537 ;
    END
    ANTENNADIFFAREA 2.4808 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.435 1.027 0.477 1.069 ;
        RECT 0.739 1.027 0.781 1.069 ;
        RECT 1.043 1.027 1.085 1.069 ;
        RECT 1.347 1.027 1.389 1.069 ;
        RECT 1.651 1.027 1.693 1.069 ;
        RECT 1.955 1.027 1.997 1.069 ;
        RECT 2.259 1.027 2.301 1.069 ;
        RECT 2.563 1.027 2.605 1.069 ;
        RECT 2.867 1.027 2.909 1.069 ;
        RECT 3.171 1.027 3.213 1.069 ;
        RECT 3.475 1.027 3.517 1.069 ;
        RECT 3.779 1.027 3.821 1.069 ;
        RECT 4.083 1.027 4.125 1.069 ;
        RECT 4.387 1.027 4.429 1.069 ;
        RECT 4.691 1.027 4.733 1.069 ;
        RECT 4.995 1.027 5.037 1.069 ;
        RECT 5.299 1.027 5.341 1.069 ;
        RECT 5.603 1.027 5.645 1.069 ;
        RECT 5.907 1.027 5.949 1.069 ;
        RECT 6.211 1.027 6.253 1.069 ;
        RECT 6.515 1.027 6.557 1.069 ;
        RECT 0.435 1.119 0.477 1.161 ;
        RECT 0.739 1.119 0.781 1.161 ;
        RECT 1.043 1.119 1.085 1.161 ;
        RECT 1.347 1.119 1.389 1.161 ;
        RECT 1.651 1.119 1.693 1.161 ;
        RECT 1.955 1.119 1.997 1.161 ;
        RECT 2.259 1.119 2.301 1.161 ;
        RECT 2.563 1.119 2.605 1.161 ;
        RECT 2.867 1.119 2.909 1.161 ;
        RECT 3.171 1.119 3.213 1.161 ;
        RECT 3.475 1.119 3.517 1.161 ;
        RECT 3.779 1.119 3.821 1.161 ;
        RECT 4.083 1.119 4.125 1.161 ;
        RECT 4.387 1.119 4.429 1.161 ;
        RECT 4.691 1.119 4.733 1.161 ;
        RECT 4.995 1.119 5.037 1.161 ;
        RECT 5.299 1.119 5.341 1.161 ;
        RECT 5.603 1.119 5.645 1.161 ;
        RECT 5.907 1.119 5.949 1.161 ;
        RECT 6.211 1.119 6.253 1.161 ;
        RECT 6.515 1.119 6.557 1.161 ;
        RECT 0.435 1.211 0.477 1.253 ;
        RECT 0.739 1.211 0.781 1.253 ;
        RECT 1.043 1.211 1.085 1.253 ;
        RECT 1.347 1.211 1.389 1.253 ;
        RECT 1.651 1.211 1.693 1.253 ;
        RECT 1.955 1.211 1.997 1.253 ;
        RECT 2.259 1.211 2.301 1.253 ;
        RECT 2.563 1.211 2.605 1.253 ;
        RECT 2.867 1.211 2.909 1.253 ;
        RECT 3.171 1.211 3.213 1.253 ;
        RECT 3.475 1.211 3.517 1.253 ;
        RECT 3.779 1.211 3.821 1.253 ;
        RECT 4.083 1.211 4.125 1.253 ;
        RECT 4.387 1.211 4.429 1.253 ;
        RECT 4.691 1.211 4.733 1.253 ;
        RECT 4.995 1.211 5.037 1.253 ;
        RECT 5.299 1.211 5.341 1.253 ;
        RECT 5.603 1.211 5.645 1.253 ;
        RECT 5.907 1.211 5.949 1.253 ;
        RECT 6.211 1.211 6.253 1.253 ;
        RECT 6.515 1.211 6.557 1.253 ;
        RECT 0.435 1.303 0.477 1.345 ;
        RECT 0.739 1.303 0.781 1.345 ;
        RECT 1.043 1.303 1.085 1.345 ;
        RECT 1.347 1.303 1.389 1.345 ;
        RECT 1.651 1.303 1.693 1.345 ;
        RECT 1.955 1.303 1.997 1.345 ;
        RECT 2.259 1.303 2.301 1.345 ;
        RECT 2.563 1.303 2.605 1.345 ;
        RECT 2.867 1.303 2.909 1.345 ;
        RECT 3.171 1.303 3.213 1.345 ;
        RECT 3.475 1.303 3.517 1.345 ;
        RECT 3.779 1.303 3.821 1.345 ;
        RECT 4.083 1.303 4.125 1.345 ;
        RECT 4.387 1.303 4.429 1.345 ;
        RECT 4.691 1.303 4.733 1.345 ;
        RECT 4.995 1.303 5.037 1.345 ;
        RECT 5.299 1.303 5.341 1.345 ;
        RECT 5.603 1.303 5.645 1.345 ;
        RECT 5.907 1.303 5.949 1.345 ;
        RECT 6.211 1.303 6.253 1.345 ;
        RECT 6.515 1.303 6.557 1.345 ;
        RECT 0.435 1.395 0.477 1.437 ;
        RECT 0.739 1.395 0.781 1.437 ;
        RECT 1.043 1.395 1.085 1.437 ;
        RECT 1.347 1.395 1.389 1.437 ;
        RECT 1.651 1.395 1.693 1.437 ;
        RECT 1.955 1.395 1.997 1.437 ;
        RECT 2.259 1.395 2.301 1.437 ;
        RECT 2.563 1.395 2.605 1.437 ;
        RECT 2.867 1.395 2.909 1.437 ;
        RECT 3.171 1.395 3.213 1.437 ;
        RECT 3.475 1.395 3.517 1.437 ;
        RECT 3.779 1.395 3.821 1.437 ;
        RECT 4.083 1.395 4.125 1.437 ;
        RECT 4.387 1.395 4.429 1.437 ;
        RECT 4.691 1.395 4.733 1.437 ;
        RECT 4.995 1.395 5.037 1.437 ;
        RECT 5.299 1.395 5.341 1.437 ;
        RECT 5.603 1.395 5.645 1.437 ;
        RECT 5.907 1.395 5.949 1.437 ;
        RECT 6.211 1.395 6.253 1.437 ;
        RECT 6.515 1.395 6.557 1.437 ;
        RECT 0.435 1.487 0.477 1.529 ;
        RECT 0.739 1.487 0.781 1.529 ;
        RECT 1.043 1.487 1.085 1.529 ;
        RECT 1.347 1.487 1.389 1.529 ;
        RECT 1.651 1.487 1.693 1.529 ;
        RECT 1.955 1.487 1.997 1.529 ;
        RECT 2.259 1.487 2.301 1.529 ;
        RECT 2.563 1.487 2.605 1.529 ;
        RECT 2.867 1.487 2.909 1.529 ;
        RECT 3.171 1.487 3.213 1.529 ;
        RECT 3.475 1.487 3.517 1.529 ;
        RECT 3.779 1.487 3.821 1.529 ;
        RECT 4.083 1.487 4.125 1.529 ;
        RECT 4.387 1.487 4.429 1.529 ;
        RECT 4.691 1.487 4.733 1.529 ;
        RECT 4.995 1.487 5.037 1.529 ;
        RECT 5.299 1.487 5.341 1.529 ;
        RECT 5.603 1.487 5.645 1.529 ;
        RECT 5.907 1.487 5.949 1.529 ;
        RECT 6.211 1.487 6.253 1.529 ;
        RECT 6.515 1.487 6.557 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
        RECT 3.095 1.651 3.137 1.693 ;
        RECT 3.247 1.651 3.289 1.693 ;
        RECT 3.399 1.651 3.441 1.693 ;
        RECT 3.551 1.651 3.593 1.693 ;
        RECT 3.703 1.651 3.745 1.693 ;
        RECT 3.855 1.651 3.897 1.693 ;
        RECT 4.007 1.651 4.049 1.693 ;
        RECT 4.159 1.651 4.201 1.693 ;
        RECT 4.311 1.651 4.353 1.693 ;
        RECT 4.463 1.651 4.505 1.693 ;
        RECT 4.615 1.651 4.657 1.693 ;
        RECT 4.767 1.651 4.809 1.693 ;
        RECT 4.919 1.651 4.961 1.693 ;
        RECT 5.071 1.651 5.113 1.693 ;
        RECT 5.223 1.651 5.265 1.693 ;
        RECT 5.375 1.651 5.417 1.693 ;
        RECT 5.527 1.651 5.569 1.693 ;
        RECT 5.679 1.651 5.721 1.693 ;
        RECT 5.831 1.651 5.873 1.693 ;
        RECT 5.983 1.651 6.025 1.693 ;
        RECT 6.135 1.651 6.177 1.693 ;
        RECT 6.287 1.651 6.329 1.693 ;
        RECT 6.439 1.651 6.481 1.693 ;
        RECT 6.591 1.651 6.633 1.693 ;
        RECT 6.743 1.651 6.785 1.693 ;
        RECT 6.895 1.651 6.937 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 6.992 1.702 ;
        RECT 3.471 0.992 3.521 1.642 ;
        RECT 3.775 0.992 3.825 1.642 ;
        RECT 4.079 0.992 4.129 1.642 ;
        RECT 4.383 0.992 4.433 1.642 ;
        RECT 4.687 0.992 4.737 1.642 ;
        RECT 4.991 0.992 5.041 1.642 ;
        RECT 5.295 0.992 5.345 1.642 ;
        RECT 5.599 0.992 5.649 1.642 ;
        RECT 5.903 0.992 5.953 1.642 ;
        RECT 6.207 0.992 6.257 1.642 ;
        RECT 6.511 0.992 6.561 1.642 ;
        RECT 0.431 0.992 0.481 1.642 ;
        RECT 0.735 0.992 0.785 1.642 ;
        RECT 1.039 0.992 1.089 1.642 ;
        RECT 1.343 0.992 1.393 1.642 ;
        RECT 1.647 0.992 1.697 1.642 ;
        RECT 1.951 0.992 2.001 1.642 ;
        RECT 2.255 0.992 2.305 1.642 ;
        RECT 2.559 0.992 2.609 1.642 ;
        RECT 2.863 0.992 2.913 1.642 ;
        RECT 3.167 0.992 3.217 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 3.399 -0.021 3.441 0.021 ;
        RECT 3.551 -0.021 3.593 0.021 ;
        RECT 3.703 -0.021 3.745 0.021 ;
        RECT 3.855 -0.021 3.897 0.021 ;
        RECT 4.007 -0.021 4.049 0.021 ;
        RECT 4.159 -0.021 4.201 0.021 ;
        RECT 4.311 -0.021 4.353 0.021 ;
        RECT 4.463 -0.021 4.505 0.021 ;
        RECT 4.615 -0.021 4.657 0.021 ;
        RECT 4.767 -0.021 4.809 0.021 ;
        RECT 4.919 -0.021 4.961 0.021 ;
        RECT 5.071 -0.021 5.113 0.021 ;
        RECT 5.223 -0.021 5.265 0.021 ;
        RECT 5.375 -0.021 5.417 0.021 ;
        RECT 5.527 -0.021 5.569 0.021 ;
        RECT 5.679 -0.021 5.721 0.021 ;
        RECT 5.831 -0.021 5.873 0.021 ;
        RECT 5.983 -0.021 6.025 0.021 ;
        RECT 6.135 -0.021 6.177 0.021 ;
        RECT 6.287 -0.021 6.329 0.021 ;
        RECT 6.439 -0.021 6.481 0.021 ;
        RECT 6.591 -0.021 6.633 0.021 ;
        RECT 6.743 -0.021 6.785 0.021 ;
        RECT 6.895 -0.021 6.937 0.021 ;
        RECT 0.435 0.149 0.477 0.191 ;
        RECT 0.739 0.149 0.781 0.191 ;
        RECT 1.043 0.149 1.085 0.191 ;
        RECT 1.347 0.149 1.389 0.191 ;
        RECT 1.651 0.149 1.693 0.191 ;
        RECT 1.955 0.149 1.997 0.191 ;
        RECT 2.259 0.149 2.301 0.191 ;
        RECT 2.563 0.149 2.605 0.191 ;
        RECT 2.867 0.149 2.909 0.191 ;
        RECT 3.171 0.149 3.213 0.191 ;
        RECT 3.475 0.149 3.517 0.191 ;
        RECT 3.779 0.149 3.821 0.191 ;
        RECT 4.083 0.149 4.125 0.191 ;
        RECT 4.387 0.149 4.429 0.191 ;
        RECT 4.691 0.149 4.733 0.191 ;
        RECT 4.995 0.149 5.037 0.191 ;
        RECT 5.299 0.149 5.341 0.191 ;
        RECT 5.603 0.149 5.645 0.191 ;
        RECT 5.907 0.149 5.949 0.191 ;
        RECT 6.211 0.149 6.253 0.191 ;
        RECT 6.515 0.149 6.557 0.191 ;
        RECT 0.435 0.241 0.477 0.283 ;
        RECT 0.739 0.241 0.781 0.283 ;
        RECT 1.043 0.241 1.085 0.283 ;
        RECT 1.347 0.241 1.389 0.283 ;
        RECT 1.651 0.241 1.693 0.283 ;
        RECT 1.955 0.241 1.997 0.283 ;
        RECT 2.259 0.241 2.301 0.283 ;
        RECT 2.563 0.241 2.605 0.283 ;
        RECT 2.867 0.241 2.909 0.283 ;
        RECT 3.171 0.241 3.213 0.283 ;
        RECT 3.475 0.241 3.517 0.283 ;
        RECT 3.779 0.241 3.821 0.283 ;
        RECT 4.083 0.241 4.125 0.283 ;
        RECT 4.387 0.241 4.429 0.283 ;
        RECT 4.691 0.241 4.733 0.283 ;
        RECT 4.995 0.241 5.037 0.283 ;
        RECT 5.299 0.241 5.341 0.283 ;
        RECT 5.603 0.241 5.645 0.283 ;
        RECT 5.907 0.241 5.949 0.283 ;
        RECT 6.211 0.241 6.253 0.283 ;
        RECT 6.515 0.241 6.557 0.283 ;
        RECT 0.435 0.333 0.477 0.375 ;
        RECT 0.739 0.333 0.781 0.375 ;
        RECT 1.043 0.333 1.085 0.375 ;
        RECT 1.347 0.333 1.389 0.375 ;
        RECT 1.651 0.333 1.693 0.375 ;
        RECT 1.955 0.333 1.997 0.375 ;
        RECT 2.259 0.333 2.301 0.375 ;
        RECT 2.563 0.333 2.605 0.375 ;
        RECT 2.867 0.333 2.909 0.375 ;
        RECT 3.171 0.333 3.213 0.375 ;
        RECT 3.475 0.333 3.517 0.375 ;
        RECT 3.779 0.333 3.821 0.375 ;
        RECT 4.083 0.333 4.125 0.375 ;
        RECT 4.387 0.333 4.429 0.375 ;
        RECT 4.691 0.333 4.733 0.375 ;
        RECT 4.995 0.333 5.037 0.375 ;
        RECT 5.299 0.333 5.341 0.375 ;
        RECT 5.603 0.333 5.645 0.375 ;
        RECT 5.907 0.333 5.949 0.375 ;
        RECT 6.211 0.333 6.253 0.375 ;
        RECT 6.515 0.333 6.557 0.375 ;
      LAYER M1 ;
        RECT 3.471 0.03 3.521 0.41 ;
        RECT 0 -0.03 6.992 0.03 ;
        RECT 3.775 0.03 3.825 0.41 ;
        RECT 4.079 0.03 4.129 0.41 ;
        RECT 4.383 0.03 4.433 0.41 ;
        RECT 4.687 0.03 4.737 0.41 ;
        RECT 4.991 0.03 5.041 0.41 ;
        RECT 5.295 0.03 5.345 0.41 ;
        RECT 5.599 0.03 5.649 0.41 ;
        RECT 5.903 0.03 5.953 0.41 ;
        RECT 6.207 0.03 6.257 0.41 ;
        RECT 6.511 0.03 6.561 0.41 ;
        RECT 0.431 0.03 0.481 0.41 ;
        RECT 0.735 0.03 0.785 0.41 ;
        RECT 1.039 0.03 1.089 0.41 ;
        RECT 1.343 0.03 1.393 0.41 ;
        RECT 1.647 0.03 1.697 0.41 ;
        RECT 1.951 0.03 2.001 0.41 ;
        RECT 2.255 0.03 2.305 0.41 ;
        RECT 2.559 0.03 2.609 0.41 ;
        RECT 2.863 0.03 2.913 0.41 ;
        RECT 3.167 0.03 3.217 0.41 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.283 1.211 0.325 1.253 ;
      RECT 0.587 1.211 0.629 1.253 ;
      RECT 0.283 1.211 0.325 1.253 ;
      RECT 0.587 1.303 0.629 1.345 ;
      RECT 0.587 0.151 0.629 0.193 ;
      RECT 0.587 1.027 0.629 1.069 ;
      RECT 1.195 0.151 1.237 0.193 ;
      RECT 1.195 1.027 1.237 1.069 ;
      RECT 1.195 0.427 1.237 0.469 ;
      RECT 1.195 0.335 1.237 0.377 ;
      RECT 1.195 1.119 1.237 1.161 ;
      RECT 1.195 1.027 1.237 1.069 ;
      RECT 0.587 0.243 0.629 0.285 ;
      RECT 0.587 1.487 0.629 1.529 ;
      RECT 0.587 0.335 0.629 0.377 ;
      RECT 1.195 0.335 1.237 0.377 ;
      RECT 1.195 1.487 1.237 1.529 ;
      RECT 1.195 0.243 1.237 0.285 ;
      RECT 1.499 1.027 1.541 1.069 ;
      RECT 1.195 1.487 1.237 1.529 ;
      RECT 1.195 1.395 1.237 1.437 ;
      RECT 1.195 0.151 1.237 0.193 ;
      RECT 0.815 0.664 0.857 0.706 ;
      RECT 0.587 0.427 0.629 0.469 ;
      RECT 1.195 1.119 1.237 1.161 ;
      RECT 1.195 1.395 1.237 1.437 ;
      RECT 1.195 1.211 1.237 1.253 ;
      RECT 0.587 1.487 0.629 1.529 ;
      RECT 1.499 1.487 1.541 1.529 ;
      RECT 1.195 1.211 1.237 1.253 ;
      RECT 1.119 0.664 1.161 0.706 ;
      RECT 1.195 1.303 1.237 1.345 ;
      RECT 0.587 0.335 0.629 0.377 ;
      RECT 6.591 0.664 6.633 0.706 ;
      RECT 5.223 0.664 5.265 0.706 ;
      RECT 4.919 0.664 4.961 0.706 ;
      RECT 5.071 0.664 5.113 0.706 ;
      RECT 4.767 0.664 4.809 0.706 ;
      RECT 4.615 0.664 4.657 0.706 ;
      RECT 4.463 0.664 4.505 0.706 ;
      RECT 4.311 0.664 4.353 0.706 ;
      RECT 5.983 0.664 6.025 0.706 ;
      RECT 6.439 0.664 6.481 0.706 ;
      RECT 6.135 0.664 6.177 0.706 ;
      RECT 6.287 0.664 6.329 0.706 ;
      RECT 5.375 0.664 5.417 0.706 ;
      RECT 5.831 0.664 5.873 0.706 ;
      RECT 5.527 0.664 5.569 0.706 ;
      RECT 0.967 0.664 1.009 0.706 ;
      RECT 1.195 1.303 1.237 1.345 ;
      RECT 1.499 1.303 1.541 1.345 ;
      RECT 1.499 1.303 1.541 1.345 ;
      RECT 1.499 1.487 1.541 1.529 ;
      RECT 1.499 1.211 1.541 1.253 ;
      RECT 1.499 1.211 1.541 1.253 ;
      RECT 1.499 1.395 1.541 1.437 ;
      RECT 1.499 1.119 1.541 1.161 ;
      RECT 1.499 1.119 1.541 1.161 ;
      RECT 1.499 1.395 1.541 1.437 ;
      RECT 1.499 1.027 1.541 1.069 ;
      RECT 0.891 1.027 0.933 1.069 ;
      RECT 0.891 1.119 0.933 1.161 ;
      RECT 0.891 1.027 0.933 1.069 ;
      RECT 0.891 1.487 0.933 1.529 ;
      RECT 0.891 1.487 0.933 1.529 ;
      RECT 0.891 1.395 0.933 1.437 ;
      RECT 0.891 1.119 0.933 1.161 ;
      RECT 0.891 1.395 0.933 1.437 ;
      RECT 0.891 1.211 0.933 1.253 ;
      RECT 0.891 1.211 0.933 1.253 ;
      RECT 0.891 1.303 0.933 1.345 ;
      RECT 0.891 1.303 0.933 1.345 ;
      RECT 0.891 0.151 0.933 0.193 ;
      RECT 0.891 0.427 0.933 0.469 ;
      RECT 0.891 0.335 0.933 0.377 ;
      RECT 0.891 0.335 0.933 0.377 ;
      RECT 0.891 0.243 0.933 0.285 ;
      RECT 0.891 0.151 0.933 0.193 ;
      RECT 1.499 0.151 1.541 0.193 ;
      RECT 1.499 0.427 1.541 0.469 ;
      RECT 1.499 0.335 1.541 0.377 ;
      RECT 1.499 0.335 1.541 0.377 ;
      RECT 1.499 0.243 1.541 0.285 ;
      RECT 1.499 0.151 1.541 0.193 ;
      RECT 1.271 0.664 1.313 0.706 ;
      RECT 1.423 0.664 1.465 0.706 ;
      RECT 1.575 0.664 1.617 0.706 ;
      RECT 0.283 1.303 0.325 1.345 ;
      RECT 0.587 1.211 0.629 1.253 ;
      RECT 0.587 1.395 0.629 1.437 ;
      RECT 0.587 1.027 0.629 1.069 ;
      RECT 0.587 1.119 0.629 1.161 ;
      RECT 0.587 0.151 0.629 0.193 ;
      RECT 0.283 0.151 0.325 0.193 ;
      RECT 0.283 1.395 0.325 1.437 ;
      RECT 0.283 1.487 0.325 1.529 ;
      RECT 0.587 1.119 0.629 1.161 ;
      RECT 0.283 0.427 0.325 0.469 ;
      RECT 5.679 0.664 5.721 0.706 ;
      RECT 0.587 1.303 0.629 1.345 ;
      RECT 0.283 0.335 0.325 0.377 ;
      RECT 0.283 0.335 0.325 0.377 ;
      RECT 0.587 1.395 0.629 1.437 ;
      RECT 3.703 0.664 3.745 0.706 ;
      RECT 4.159 0.664 4.201 0.706 ;
      RECT 3.855 0.664 3.897 0.706 ;
      RECT 4.007 0.664 4.049 0.706 ;
      RECT 0.283 0.243 0.325 0.285 ;
      RECT 0.283 1.395 0.325 1.437 ;
      RECT 0.283 1.027 0.325 1.069 ;
      RECT 3.095 0.664 3.137 0.706 ;
      RECT 3.551 0.664 3.593 0.706 ;
      RECT 3.247 0.664 3.289 0.706 ;
      RECT 3.399 0.664 3.441 0.706 ;
      RECT 0.283 1.119 0.325 1.161 ;
      RECT 0.283 1.303 0.325 1.345 ;
      RECT 1.879 0.664 1.921 0.706 ;
      RECT 2.031 0.664 2.073 0.706 ;
      RECT 0.283 1.487 0.325 1.529 ;
      RECT 0.283 1.027 0.325 1.069 ;
      RECT 0.283 1.119 0.325 1.161 ;
      RECT 2.639 0.664 2.681 0.706 ;
      RECT 2.791 0.664 2.833 0.706 ;
      RECT 2.487 0.664 2.529 0.706 ;
      RECT 0.283 0.151 0.325 0.193 ;
      RECT 2.335 0.664 2.377 0.706 ;
      RECT 2.183 0.664 2.225 0.706 ;
      RECT 2.943 0.664 2.985 0.706 ;
    LAYER M1 ;
      RECT 1.702 0.66 6.668 0.71 ;
      RECT 0.887 0.942 0.937 1.564 ;
      RECT 0.887 0.116 0.937 0.537 ;
      RECT 1.191 0.942 1.241 1.564 ;
      RECT 1.191 0.116 1.241 0.537 ;
      RECT 1.495 0.942 1.545 1.564 ;
      RECT 1.495 0.116 1.545 0.537 ;
      RECT 0.887 0.537 1.749 0.587 ;
      RECT 1.702 0.71 1.752 0.818 ;
      RECT 1.699 0.874 1.749 0.892 ;
      RECT 1.699 0.818 1.752 0.874 ;
      RECT 1.699 0.587 1.749 0.605 ;
      RECT 1.702 0.631 1.752 0.66 ;
      RECT 1.699 0.605 1.752 0.631 ;
      RECT 0.887 0.892 1.749 0.942 ;
      RECT 0.639 0.66 1.652 0.71 ;
      RECT 0.279 0.116 0.329 0.537 ;
      RECT 0.279 0.942 0.329 1.564 ;
      RECT 0.583 0.942 0.633 1.564 ;
      RECT 0.279 0.537 0.689 0.587 ;
      RECT 0.639 0.587 0.689 0.66 ;
      RECT 0.583 0.116 0.633 0.537 ;
      RECT 0.639 0.71 0.689 0.892 ;
      RECT 0.279 0.892 0.689 0.942 ;
    LAYER PO ;
      RECT 1.885 0.069 1.915 1.606 ;
      RECT 2.341 0.069 2.371 1.606 ;
      RECT 2.189 0.069 2.219 1.606 ;
      RECT 2.037 0.069 2.067 1.606 ;
      RECT 0.061 0.071 0.091 1.606 ;
      RECT 0.669 0.069 0.699 1.606 ;
      RECT 0.517 0.069 0.547 1.606 ;
      RECT 1.125 0.069 1.155 1.606 ;
      RECT 1.277 0.069 1.307 1.606 ;
      RECT 1.429 0.069 1.459 1.606 ;
      RECT 0.973 0.069 1.003 1.606 ;
      RECT 0.821 0.069 0.851 1.606 ;
      RECT 1.581 0.069 1.611 1.606 ;
      RECT 0.213 0.071 0.243 1.606 ;
      RECT 0.365 0.069 0.395 1.606 ;
      RECT 6.901 0.069 6.931 1.606 ;
      RECT 6.749 0.069 6.779 1.606 ;
      RECT 6.597 0.069 6.627 1.606 ;
      RECT 6.445 0.069 6.475 1.606 ;
      RECT 6.141 0.069 6.171 1.606 ;
      RECT 6.293 0.069 6.323 1.606 ;
      RECT 5.837 0.069 5.867 1.606 ;
      RECT 5.989 0.069 6.019 1.606 ;
      RECT 5.685 0.069 5.715 1.606 ;
      RECT 5.533 0.069 5.563 1.606 ;
      RECT 5.381 0.069 5.411 1.606 ;
      RECT 5.229 0.069 5.259 1.606 ;
      RECT 4.925 0.069 4.955 1.606 ;
      RECT 5.077 0.069 5.107 1.606 ;
      RECT 4.317 0.069 4.347 1.606 ;
      RECT 4.469 0.069 4.499 1.606 ;
      RECT 4.165 0.069 4.195 1.606 ;
      RECT 4.621 0.069 4.651 1.606 ;
      RECT 4.773 0.069 4.803 1.606 ;
      RECT 2.949 0.069 2.979 1.606 ;
      RECT 3.101 0.069 3.131 1.606 ;
      RECT 3.253 0.069 3.283 1.606 ;
      RECT 3.861 0.069 3.891 1.606 ;
      RECT 3.709 0.069 3.739 1.606 ;
      RECT 3.557 0.069 3.587 1.606 ;
      RECT 3.405 0.069 3.435 1.606 ;
      RECT 4.013 0.069 4.043 1.606 ;
      RECT 2.797 0.069 2.827 1.606 ;
      RECT 2.645 0.069 2.675 1.606 ;
      RECT 2.493 0.069 2.523 1.606 ;
      RECT 1.733 0.069 1.763 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 7.107 1.773 ;
  END
END IBUFFX32_RVT

MACRO IBUFFX8_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.684 0.401 0.726 ;
      LAYER M1 ;
        RECT 0.249 0.73 0.362 0.815 ;
        RECT 0.249 0.68 0.436 0.73 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.043 0.151 1.085 0.193 ;
        RECT 1.347 0.151 1.389 0.193 ;
        RECT 1.651 0.151 1.693 0.193 ;
        RECT 1.955 0.151 1.997 0.193 ;
        RECT 2.259 0.152 2.301 0.194 ;
        RECT 1.043 0.243 1.085 0.285 ;
        RECT 1.347 0.243 1.389 0.285 ;
        RECT 1.651 0.243 1.693 0.285 ;
        RECT 1.955 0.243 1.997 0.285 ;
        RECT 2.259 0.244 2.301 0.286 ;
        RECT 1.043 0.335 1.085 0.377 ;
        RECT 1.347 0.335 1.389 0.377 ;
        RECT 1.651 0.335 1.693 0.377 ;
        RECT 1.955 0.335 1.997 0.377 ;
        RECT 2.259 0.336 2.301 0.378 ;
        RECT 1.043 0.427 1.085 0.469 ;
        RECT 1.347 0.427 1.389 0.469 ;
        RECT 1.651 0.427 1.693 0.469 ;
        RECT 1.955 0.427 1.997 0.469 ;
        RECT 2.259 0.428 2.301 0.47 ;
        RECT 1.043 1.027 1.085 1.069 ;
        RECT 1.347 1.027 1.389 1.069 ;
        RECT 1.651 1.027 1.693 1.069 ;
        RECT 1.955 1.027 1.997 1.069 ;
        RECT 2.259 1.028 2.301 1.07 ;
        RECT 1.043 1.119 1.085 1.161 ;
        RECT 1.347 1.119 1.389 1.161 ;
        RECT 1.651 1.119 1.693 1.161 ;
        RECT 1.955 1.119 1.997 1.161 ;
        RECT 2.259 1.12 2.301 1.162 ;
        RECT 1.043 1.211 1.085 1.253 ;
        RECT 1.347 1.211 1.389 1.253 ;
        RECT 1.651 1.211 1.693 1.253 ;
        RECT 1.955 1.211 1.997 1.253 ;
        RECT 2.259 1.212 2.301 1.254 ;
        RECT 1.043 1.303 1.085 1.345 ;
        RECT 1.347 1.303 1.389 1.345 ;
        RECT 1.651 1.303 1.693 1.345 ;
        RECT 1.955 1.303 1.997 1.345 ;
        RECT 2.259 1.304 2.301 1.346 ;
        RECT 1.043 1.395 1.085 1.437 ;
        RECT 1.347 1.395 1.389 1.437 ;
        RECT 1.651 1.395 1.693 1.437 ;
        RECT 1.955 1.395 1.997 1.437 ;
        RECT 2.259 1.396 2.301 1.438 ;
        RECT 1.043 1.487 1.085 1.529 ;
        RECT 1.347 1.487 1.389 1.529 ;
        RECT 1.651 1.487 1.693 1.529 ;
        RECT 1.955 1.487 1.997 1.529 ;
        RECT 2.259 1.488 2.301 1.53 ;
      LAYER M1 ;
        RECT 2.255 0.942 2.305 1.565 ;
        RECT 1.039 0.942 1.089 1.564 ;
        RECT 1.343 0.942 1.393 1.564 ;
        RECT 1.647 0.942 1.697 1.564 ;
        RECT 1.951 0.942 2.001 1.564 ;
        RECT 1.039 0.892 2.361 0.942 ;
        RECT 2.311 0.663 2.361 0.892 ;
        RECT 2.311 0.587 2.487 0.663 ;
        RECT 1.039 0.537 2.487 0.587 ;
        RECT 1.039 0.116 1.089 0.537 ;
        RECT 1.343 0.116 1.393 0.537 ;
        RECT 1.647 0.116 1.697 0.537 ;
        RECT 1.951 0.116 2.001 0.537 ;
        RECT 2.255 0.117 2.305 0.537 ;
    END
    ANTENNADIFFAREA 0.6952 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.435 1.027 0.477 1.069 ;
        RECT 0.739 1.027 0.781 1.069 ;
        RECT 1.195 1.027 1.237 1.069 ;
        RECT 1.499 1.027 1.541 1.069 ;
        RECT 1.803 1.027 1.845 1.069 ;
        RECT 2.107 1.027 2.149 1.069 ;
        RECT 0.435 1.119 0.477 1.161 ;
        RECT 0.739 1.119 0.781 1.161 ;
        RECT 1.195 1.119 1.237 1.161 ;
        RECT 1.499 1.119 1.541 1.161 ;
        RECT 1.803 1.119 1.845 1.161 ;
        RECT 2.107 1.119 2.149 1.161 ;
        RECT 0.435 1.211 0.477 1.253 ;
        RECT 0.739 1.211 0.781 1.253 ;
        RECT 1.195 1.211 1.237 1.253 ;
        RECT 1.499 1.211 1.541 1.253 ;
        RECT 1.803 1.211 1.845 1.253 ;
        RECT 2.107 1.211 2.149 1.253 ;
        RECT 0.739 1.303 0.781 1.345 ;
        RECT 1.195 1.303 1.237 1.345 ;
        RECT 1.499 1.303 1.541 1.345 ;
        RECT 1.803 1.303 1.845 1.345 ;
        RECT 2.107 1.303 2.149 1.345 ;
        RECT 0.739 1.395 0.781 1.437 ;
        RECT 1.195 1.395 1.237 1.437 ;
        RECT 1.499 1.395 1.541 1.437 ;
        RECT 1.803 1.395 1.845 1.437 ;
        RECT 2.107 1.395 2.149 1.437 ;
        RECT 0.739 1.487 0.781 1.529 ;
        RECT 1.195 1.487 1.237 1.529 ;
        RECT 1.499 1.487 1.541 1.529 ;
        RECT 1.803 1.487 1.845 1.529 ;
        RECT 2.107 1.487 2.149 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 2.584 1.702 ;
        RECT 0.431 0.992 0.481 1.642 ;
        RECT 0.735 0.992 0.785 1.642 ;
        RECT 1.191 0.992 1.241 1.642 ;
        RECT 1.495 0.992 1.545 1.642 ;
        RECT 1.799 0.992 1.849 1.642 ;
        RECT 2.103 0.992 2.153 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 0.739 0.149 0.781 0.191 ;
        RECT 1.195 0.149 1.237 0.191 ;
        RECT 1.499 0.149 1.541 0.191 ;
        RECT 1.803 0.149 1.845 0.191 ;
        RECT 2.107 0.149 2.149 0.191 ;
        RECT 0.739 0.241 0.781 0.283 ;
        RECT 1.195 0.241 1.237 0.283 ;
        RECT 1.499 0.241 1.541 0.283 ;
        RECT 1.803 0.241 1.845 0.283 ;
        RECT 2.107 0.241 2.149 0.283 ;
        RECT 0.435 0.318 0.477 0.36 ;
        RECT 0.739 0.333 0.781 0.375 ;
        RECT 1.195 0.333 1.237 0.375 ;
        RECT 1.499 0.333 1.541 0.375 ;
        RECT 1.803 0.333 1.845 0.375 ;
        RECT 2.107 0.333 2.149 0.375 ;
        RECT 0.435 0.41 0.477 0.452 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.487 ;
        RECT 0.735 0.03 0.785 0.41 ;
        RECT 1.191 0.03 1.241 0.41 ;
        RECT 1.495 0.03 1.545 0.41 ;
        RECT 1.799 0.03 1.849 0.41 ;
        RECT 2.103 0.03 2.153 0.41 ;
        RECT 0 -0.03 2.584 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.587 1.487 0.629 1.529 ;
      RECT 0.283 1.211 0.325 1.253 ;
      RECT 0.283 0.325 0.325 0.367 ;
      RECT 0.891 0.151 0.933 0.193 ;
      RECT 0.891 1.027 0.933 1.069 ;
      RECT 0.891 0.427 0.933 0.469 ;
      RECT 0.891 0.335 0.933 0.377 ;
      RECT 0.891 1.119 0.933 1.161 ;
      RECT 0.283 1.211 0.325 1.253 ;
      RECT 0.891 1.027 0.933 1.069 ;
      RECT 0.283 1.119 0.325 1.161 ;
      RECT 0.283 1.119 0.325 1.161 ;
      RECT 0.283 1.027 0.325 1.069 ;
      RECT 0.891 0.335 0.933 0.377 ;
      RECT 0.891 1.487 0.933 1.529 ;
      RECT 0.891 0.243 0.933 0.285 ;
      RECT 0.891 1.487 0.933 1.529 ;
      RECT 0.891 1.395 0.933 1.437 ;
      RECT 0.891 0.151 0.933 0.193 ;
      RECT 0.283 1.027 0.325 1.069 ;
      RECT 0.891 1.119 0.933 1.161 ;
      RECT 0.891 1.395 0.933 1.437 ;
      RECT 0.891 1.211 0.933 1.253 ;
      RECT 0.283 0.935 0.325 0.977 ;
      RECT 0.283 0.509 0.325 0.551 ;
      RECT 0.283 0.935 0.325 0.977 ;
      RECT 2.183 0.664 2.225 0.706 ;
      RECT 0.587 1.027 0.629 1.069 ;
      RECT 0.587 1.119 0.629 1.161 ;
      RECT 0.587 1.487 0.629 1.529 ;
      RECT 0.587 1.395 0.629 1.437 ;
      RECT 0.587 1.119 0.629 1.161 ;
      RECT 0.587 1.395 0.629 1.437 ;
      RECT 0.891 1.303 0.933 1.345 ;
      RECT 0.815 0.664 0.857 0.706 ;
      RECT 0.891 1.211 0.933 1.253 ;
      RECT 0.283 0.417 0.325 0.459 ;
      RECT 1.879 0.664 1.921 0.706 ;
      RECT 2.031 0.664 2.073 0.706 ;
      RECT 1.727 0.664 1.769 0.706 ;
      RECT 1.575 0.664 1.617 0.706 ;
      RECT 1.423 0.664 1.465 0.706 ;
      RECT 0.587 1.211 0.629 1.253 ;
      RECT 0.587 0.427 0.629 0.469 ;
      RECT 0.587 0.151 0.629 0.193 ;
      RECT 0.587 1.303 0.629 1.345 ;
      RECT 0.587 1.303 0.629 1.345 ;
      RECT 0.587 1.027 0.629 1.069 ;
      RECT 0.587 0.335 0.629 0.377 ;
      RECT 1.119 0.664 1.161 0.706 ;
      RECT 1.271 0.664 1.313 0.706 ;
      RECT 0.587 0.335 0.629 0.377 ;
      RECT 0.587 1.211 0.629 1.253 ;
      RECT 0.587 0.151 0.629 0.193 ;
      RECT 0.587 0.243 0.629 0.285 ;
      RECT 0.663 0.664 0.705 0.706 ;
      RECT 0.283 0.417 0.325 0.459 ;
      RECT 0.891 1.303 0.933 1.345 ;
    LAYER M1 ;
      RECT 0.943 0.66 2.26 0.71 ;
      RECT 0.583 0.116 0.633 0.537 ;
      RECT 0.583 0.942 0.633 1.564 ;
      RECT 0.939 0.85 0.993 0.87 ;
      RECT 0.943 0.71 0.993 0.85 ;
      RECT 0.583 0.537 0.989 0.587 ;
      RECT 0.887 0.116 0.937 0.537 ;
      RECT 0.939 0.87 0.989 0.892 ;
      RECT 0.939 0.587 0.989 0.609 ;
      RECT 0.943 0.642 0.993 0.66 ;
      RECT 0.939 0.609 0.993 0.642 ;
      RECT 0.887 0.942 0.937 1.564 ;
      RECT 0.583 0.892 0.989 0.942 ;
      RECT 0.487 0.66 0.892 0.71 ;
      RECT 0.279 0.942 0.329 1.288 ;
      RECT 0.279 0.305 0.329 0.537 ;
      RECT 0.279 0.537 0.533 0.587 ;
      RECT 0.279 0.892 0.533 0.942 ;
      RECT 0.483 0.609 0.537 0.649 ;
      RECT 0.487 0.649 0.537 0.66 ;
      RECT 0.483 0.587 0.533 0.609 ;
      RECT 0.487 0.71 0.537 0.811 ;
      RECT 0.483 0.87 0.533 0.892 ;
      RECT 0.483 0.811 0.537 0.87 ;
    LAYER PO ;
      RECT 0.061 0.071 0.091 1.606 ;
      RECT 0.365 0.069 0.395 1.606 ;
      RECT 0.213 0.071 0.243 1.606 ;
      RECT 0.821 0.069 0.851 1.606 ;
      RECT 2.189 0.069 2.219 1.606 ;
      RECT 2.341 0.069 2.371 1.606 ;
      RECT 2.493 0.069 2.523 1.606 ;
      RECT 0.517 0.071 0.547 1.606 ;
      RECT 0.669 0.069 0.699 1.606 ;
      RECT 2.037 0.069 2.067 1.606 ;
      RECT 1.885 0.069 1.915 1.606 ;
      RECT 1.733 0.069 1.763 1.606 ;
      RECT 0.973 0.069 1.003 1.606 ;
      RECT 1.125 0.069 1.155 1.606 ;
      RECT 1.581 0.069 1.611 1.606 ;
      RECT 1.429 0.069 1.459 1.606 ;
      RECT 1.277 0.069 1.307 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 2.699 1.773 ;
  END
END IBUFFX8_RVT

MACRO INVX16_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.04 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.664 0.401 0.706 ;
        RECT 0.511 0.664 0.553 0.706 ;
        RECT 0.663 0.664 0.705 0.706 ;
        RECT 0.815 0.664 0.857 0.706 ;
        RECT 0.967 0.664 1.009 0.706 ;
        RECT 1.119 0.664 1.161 0.706 ;
        RECT 1.271 0.664 1.313 0.706 ;
        RECT 1.423 0.664 1.465 0.706 ;
        RECT 1.575 0.664 1.617 0.706 ;
        RECT 1.727 0.664 1.769 0.706 ;
        RECT 1.879 0.664 1.921 0.706 ;
        RECT 2.031 0.664 2.073 0.706 ;
        RECT 2.183 0.664 2.225 0.706 ;
        RECT 2.335 0.664 2.377 0.706 ;
        RECT 2.487 0.664 2.529 0.706 ;
        RECT 2.639 0.664 2.681 0.706 ;
      LAYER M1 ;
        RECT 0.249 0.71 0.362 0.815 ;
        RECT 0.249 0.66 2.716 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5856 ;
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.283 0.151 0.325 0.193 ;
        RECT 0.587 0.151 0.629 0.193 ;
        RECT 0.891 0.151 0.933 0.193 ;
        RECT 1.195 0.151 1.237 0.193 ;
        RECT 1.803 0.151 1.845 0.193 ;
        RECT 2.107 0.151 2.149 0.193 ;
        RECT 2.411 0.151 2.453 0.193 ;
        RECT 2.715 0.151 2.757 0.193 ;
        RECT 1.499 0.152 1.541 0.194 ;
        RECT 0.283 0.243 0.325 0.285 ;
        RECT 0.587 0.243 0.629 0.285 ;
        RECT 0.891 0.243 0.933 0.285 ;
        RECT 1.195 0.243 1.237 0.285 ;
        RECT 1.803 0.243 1.845 0.285 ;
        RECT 2.107 0.243 2.149 0.285 ;
        RECT 2.411 0.243 2.453 0.285 ;
        RECT 2.715 0.243 2.757 0.285 ;
        RECT 1.499 0.244 1.541 0.286 ;
        RECT 0.283 0.335 0.325 0.377 ;
        RECT 0.587 0.335 0.629 0.377 ;
        RECT 0.891 0.335 0.933 0.377 ;
        RECT 1.195 0.335 1.237 0.377 ;
        RECT 1.803 0.335 1.845 0.377 ;
        RECT 2.107 0.335 2.149 0.377 ;
        RECT 2.411 0.335 2.453 0.377 ;
        RECT 2.715 0.335 2.757 0.377 ;
        RECT 1.499 0.336 1.541 0.378 ;
        RECT 0.283 0.427 0.325 0.469 ;
        RECT 0.587 0.427 0.629 0.469 ;
        RECT 0.891 0.427 0.933 0.469 ;
        RECT 1.195 0.427 1.237 0.469 ;
        RECT 1.803 0.427 1.845 0.469 ;
        RECT 2.107 0.427 2.149 0.469 ;
        RECT 2.411 0.427 2.453 0.469 ;
        RECT 2.715 0.427 2.757 0.469 ;
        RECT 1.499 0.428 1.541 0.47 ;
        RECT 0.283 1.027 0.325 1.069 ;
        RECT 0.587 1.027 0.629 1.069 ;
        RECT 0.891 1.027 0.933 1.069 ;
        RECT 1.195 1.027 1.237 1.069 ;
        RECT 1.803 1.027 1.845 1.069 ;
        RECT 2.107 1.027 2.149 1.069 ;
        RECT 2.411 1.027 2.453 1.069 ;
        RECT 2.715 1.027 2.757 1.069 ;
        RECT 1.499 1.028 1.541 1.07 ;
        RECT 0.283 1.119 0.325 1.161 ;
        RECT 0.587 1.119 0.629 1.161 ;
        RECT 0.891 1.119 0.933 1.161 ;
        RECT 1.195 1.119 1.237 1.161 ;
        RECT 1.803 1.119 1.845 1.161 ;
        RECT 2.107 1.119 2.149 1.161 ;
        RECT 2.411 1.119 2.453 1.161 ;
        RECT 2.715 1.119 2.757 1.161 ;
        RECT 1.499 1.12 1.541 1.162 ;
        RECT 0.283 1.211 0.325 1.253 ;
        RECT 0.587 1.211 0.629 1.253 ;
        RECT 0.891 1.211 0.933 1.253 ;
        RECT 1.195 1.211 1.237 1.253 ;
        RECT 1.803 1.211 1.845 1.253 ;
        RECT 2.107 1.211 2.149 1.253 ;
        RECT 2.411 1.211 2.453 1.253 ;
        RECT 2.715 1.211 2.757 1.253 ;
        RECT 1.499 1.212 1.541 1.254 ;
        RECT 0.283 1.303 0.325 1.345 ;
        RECT 0.587 1.303 0.629 1.345 ;
        RECT 0.891 1.303 0.933 1.345 ;
        RECT 1.195 1.303 1.237 1.345 ;
        RECT 1.803 1.303 1.845 1.345 ;
        RECT 2.107 1.303 2.149 1.345 ;
        RECT 2.411 1.303 2.453 1.345 ;
        RECT 2.715 1.303 2.757 1.345 ;
        RECT 1.499 1.304 1.541 1.346 ;
        RECT 0.283 1.395 0.325 1.437 ;
        RECT 0.587 1.395 0.629 1.437 ;
        RECT 0.891 1.395 0.933 1.437 ;
        RECT 1.195 1.395 1.237 1.437 ;
        RECT 1.803 1.395 1.845 1.437 ;
        RECT 2.107 1.395 2.149 1.437 ;
        RECT 2.411 1.395 2.453 1.437 ;
        RECT 2.715 1.395 2.757 1.437 ;
        RECT 1.499 1.396 1.541 1.438 ;
        RECT 0.283 1.487 0.325 1.529 ;
        RECT 0.587 1.487 0.629 1.529 ;
        RECT 0.891 1.487 0.933 1.529 ;
        RECT 1.195 1.487 1.237 1.529 ;
        RECT 1.803 1.487 1.845 1.529 ;
        RECT 2.107 1.487 2.149 1.529 ;
        RECT 2.411 1.487 2.453 1.529 ;
        RECT 2.715 1.487 2.757 1.529 ;
        RECT 1.499 1.488 1.541 1.53 ;
      LAYER M1 ;
        RECT 1.495 0.942 1.545 1.565 ;
        RECT 0.279 0.942 0.329 1.564 ;
        RECT 0.583 0.942 0.633 1.564 ;
        RECT 0.887 0.942 0.937 1.564 ;
        RECT 1.191 0.942 1.241 1.564 ;
        RECT 1.799 0.942 1.849 1.564 ;
        RECT 2.103 0.942 2.153 1.564 ;
        RECT 2.407 0.942 2.457 1.564 ;
        RECT 2.711 0.942 2.761 1.564 ;
        RECT 0.279 0.892 2.82 0.942 ;
        RECT 2.77 0.663 2.82 0.892 ;
        RECT 2.77 0.587 2.943 0.663 ;
        RECT 0.279 0.537 2.943 0.587 ;
        RECT 0.279 0.116 0.329 0.537 ;
        RECT 0.583 0.116 0.633 0.537 ;
        RECT 0.887 0.116 0.937 0.537 ;
        RECT 1.191 0.116 1.241 0.537 ;
        RECT 1.495 0.117 1.545 0.537 ;
        RECT 1.799 0.116 1.849 0.537 ;
        RECT 2.103 0.116 2.153 0.537 ;
        RECT 2.407 0.116 2.457 0.537 ;
        RECT 2.711 0.116 2.761 0.537 ;
    END
    ANTENNADIFFAREA 1.2904 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.435 1.027 0.477 1.069 ;
        RECT 0.739 1.027 0.781 1.069 ;
        RECT 1.043 1.027 1.085 1.069 ;
        RECT 1.347 1.027 1.389 1.069 ;
        RECT 1.651 1.027 1.693 1.069 ;
        RECT 1.955 1.027 1.997 1.069 ;
        RECT 2.259 1.027 2.301 1.069 ;
        RECT 2.563 1.027 2.605 1.069 ;
        RECT 0.435 1.119 0.477 1.161 ;
        RECT 0.739 1.119 0.781 1.161 ;
        RECT 1.043 1.119 1.085 1.161 ;
        RECT 1.347 1.119 1.389 1.161 ;
        RECT 1.651 1.119 1.693 1.161 ;
        RECT 1.955 1.119 1.997 1.161 ;
        RECT 2.259 1.119 2.301 1.161 ;
        RECT 2.563 1.119 2.605 1.161 ;
        RECT 0.435 1.211 0.477 1.253 ;
        RECT 0.739 1.211 0.781 1.253 ;
        RECT 1.043 1.211 1.085 1.253 ;
        RECT 1.347 1.211 1.389 1.253 ;
        RECT 1.651 1.211 1.693 1.253 ;
        RECT 1.955 1.211 1.997 1.253 ;
        RECT 2.259 1.211 2.301 1.253 ;
        RECT 2.563 1.211 2.605 1.253 ;
        RECT 0.435 1.303 0.477 1.345 ;
        RECT 0.739 1.303 0.781 1.345 ;
        RECT 1.043 1.303 1.085 1.345 ;
        RECT 1.347 1.303 1.389 1.345 ;
        RECT 1.651 1.303 1.693 1.345 ;
        RECT 1.955 1.303 1.997 1.345 ;
        RECT 2.259 1.303 2.301 1.345 ;
        RECT 2.563 1.303 2.605 1.345 ;
        RECT 0.435 1.395 0.477 1.437 ;
        RECT 0.739 1.395 0.781 1.437 ;
        RECT 1.043 1.395 1.085 1.437 ;
        RECT 1.347 1.395 1.389 1.437 ;
        RECT 1.651 1.395 1.693 1.437 ;
        RECT 1.955 1.395 1.997 1.437 ;
        RECT 2.259 1.395 2.301 1.437 ;
        RECT 2.563 1.395 2.605 1.437 ;
        RECT 0.435 1.487 0.477 1.529 ;
        RECT 0.739 1.487 0.781 1.529 ;
        RECT 1.043 1.487 1.085 1.529 ;
        RECT 1.347 1.487 1.389 1.529 ;
        RECT 1.651 1.487 1.693 1.529 ;
        RECT 1.955 1.487 1.997 1.529 ;
        RECT 2.259 1.487 2.301 1.529 ;
        RECT 2.563 1.487 2.605 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 3.04 1.702 ;
        RECT 0.431 0.992 0.481 1.642 ;
        RECT 0.735 0.992 0.785 1.642 ;
        RECT 1.039 0.992 1.089 1.642 ;
        RECT 1.343 0.992 1.393 1.642 ;
        RECT 1.647 0.992 1.697 1.642 ;
        RECT 1.951 0.992 2.001 1.642 ;
        RECT 2.255 0.992 2.305 1.642 ;
        RECT 2.559 0.992 2.609 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 0.435 0.149 0.477 0.191 ;
        RECT 0.739 0.149 0.781 0.191 ;
        RECT 1.043 0.149 1.085 0.191 ;
        RECT 1.347 0.149 1.389 0.191 ;
        RECT 1.651 0.149 1.693 0.191 ;
        RECT 1.955 0.149 1.997 0.191 ;
        RECT 2.259 0.149 2.301 0.191 ;
        RECT 2.563 0.149 2.605 0.191 ;
        RECT 0.435 0.241 0.477 0.283 ;
        RECT 0.739 0.241 0.781 0.283 ;
        RECT 1.043 0.241 1.085 0.283 ;
        RECT 1.347 0.241 1.389 0.283 ;
        RECT 1.651 0.241 1.693 0.283 ;
        RECT 1.955 0.241 1.997 0.283 ;
        RECT 2.259 0.241 2.301 0.283 ;
        RECT 2.563 0.241 2.605 0.283 ;
        RECT 0.435 0.333 0.477 0.375 ;
        RECT 0.739 0.333 0.781 0.375 ;
        RECT 1.043 0.333 1.085 0.375 ;
        RECT 1.347 0.333 1.389 0.375 ;
        RECT 1.651 0.333 1.693 0.375 ;
        RECT 1.955 0.333 1.997 0.375 ;
        RECT 2.259 0.333 2.301 0.375 ;
        RECT 2.563 0.333 2.605 0.375 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.41 ;
        RECT 0.735 0.03 0.785 0.41 ;
        RECT 1.039 0.03 1.089 0.41 ;
        RECT 1.343 0.03 1.393 0.41 ;
        RECT 1.647 0.03 1.697 0.41 ;
        RECT 1.951 0.03 2.001 0.41 ;
        RECT 2.255 0.03 2.305 0.41 ;
        RECT 2.559 0.03 2.609 0.41 ;
        RECT 0 -0.03 3.04 0.03 ;
    END
  END VSS
  OBS
    LAYER PO ;
      RECT 2.797 0.069 2.827 1.606 ;
      RECT 2.949 0.069 2.979 1.606 ;
      RECT 2.645 0.069 2.675 1.606 ;
      RECT 1.429 0.069 1.459 1.606 ;
      RECT 1.581 0.069 1.611 1.606 ;
      RECT 1.733 0.069 1.763 1.606 ;
      RECT 2.341 0.069 2.371 1.606 ;
      RECT 2.189 0.069 2.219 1.606 ;
      RECT 2.037 0.069 2.067 1.606 ;
      RECT 1.885 0.069 1.915 1.606 ;
      RECT 2.493 0.069 2.523 1.606 ;
      RECT 1.277 0.069 1.307 1.606 ;
      RECT 1.125 0.069 1.155 1.606 ;
      RECT 0.973 0.069 1.003 1.606 ;
      RECT 0.213 0.069 0.243 1.606 ;
      RECT 0.365 0.069 0.395 1.606 ;
      RECT 0.821 0.069 0.851 1.606 ;
      RECT 0.669 0.069 0.699 1.606 ;
      RECT 0.517 0.069 0.547 1.606 ;
      RECT 0.061 0.069 0.091 1.606 ;
    LAYER NWELL ;
      RECT -0.115 0.679 3.155 1.773 ;
  END
END INVX16_RVT

MACRO MUX21X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.615 0.401 0.657 ;
      LAYER M1 ;
        RECT 0.355 0.663 0.405 0.692 ;
        RECT 0.23 0.553 0.415 0.663 ;
        RECT 0.355 0.499 0.405 0.553 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.271 0.891 1.313 0.933 ;
      LAYER M1 ;
        RECT 1.251 0.857 1.423 0.967 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 ;
  END A2
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.119 0.634 1.161 0.676 ;
        RECT 0.815 0.733 0.857 0.775 ;
        RECT 0.511 0.967 0.553 1.009 ;
      LAYER M1 ;
        RECT 0.507 0.755 0.557 1.029 ;
        RECT 0.811 0.755 0.967 0.815 ;
        RECT 0.507 0.705 0.967 0.755 ;
        RECT 0.507 0.663 0.557 0.705 ;
        RECT 0.917 0.664 0.967 0.705 ;
        RECT 1.115 0.664 1.165 0.696 ;
        RECT 0.917 0.614 1.165 0.664 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.651 0.152 1.693 0.194 ;
        RECT 1.651 0.244 1.693 0.286 ;
        RECT 1.651 0.336 1.693 0.378 ;
        RECT 1.651 0.428 1.693 0.47 ;
        RECT 1.651 0.931 1.693 0.973 ;
        RECT 1.651 1.023 1.693 1.065 ;
        RECT 1.651 1.115 1.693 1.157 ;
        RECT 1.651 1.207 1.693 1.249 ;
        RECT 1.651 1.299 1.693 1.341 ;
        RECT 1.651 1.391 1.693 1.433 ;
        RECT 1.651 1.483 1.693 1.525 ;
      LAYER M1 ;
        RECT 1.647 0.885 1.697 1.545 ;
        RECT 1.647 0.835 1.959 0.885 ;
        RECT 1.909 0.815 1.959 0.835 ;
        RECT 1.909 0.705 2.038 0.815 ;
        RECT 1.909 0.498 1.959 0.705 ;
        RECT 1.647 0.448 1.959 0.498 ;
        RECT 1.647 0.132 1.697 0.448 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.803 1.023 1.845 1.065 ;
        RECT 1.803 1.115 1.845 1.157 ;
        RECT 1.803 1.207 1.845 1.249 ;
        RECT 1.499 1.299 1.541 1.341 ;
        RECT 1.803 1.299 1.845 1.341 ;
        RECT 0.587 1.312 0.629 1.354 ;
        RECT 0.891 1.313 0.933 1.355 ;
        RECT 1.043 1.313 1.085 1.355 ;
        RECT 1.499 1.391 1.541 1.433 ;
        RECT 1.803 1.391 1.845 1.433 ;
        RECT 0.587 1.404 0.629 1.446 ;
        RECT 0.891 1.405 0.933 1.447 ;
        RECT 1.043 1.405 1.085 1.447 ;
        RECT 1.499 1.483 1.541 1.525 ;
        RECT 1.803 1.483 1.845 1.525 ;
        RECT 0.587 1.496 0.629 1.538 ;
        RECT 0.891 1.497 0.933 1.539 ;
        RECT 1.043 1.497 1.085 1.539 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 2.128 1.702 ;
        RECT 0.583 1.292 0.633 1.642 ;
        RECT 0.887 1.292 0.937 1.642 ;
        RECT 1.039 1.292 1.089 1.642 ;
        RECT 1.495 1.279 1.545 1.642 ;
        RECT 1.799 1.003 1.849 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 0.587 0.141 0.629 0.183 ;
        RECT 0.891 0.142 0.933 0.184 ;
        RECT 1.043 0.142 1.085 0.184 ;
        RECT 1.499 0.16 1.541 0.202 ;
        RECT 1.803 0.16 1.845 0.202 ;
        RECT 0.587 0.233 0.629 0.275 ;
        RECT 0.891 0.234 0.933 0.276 ;
        RECT 1.043 0.234 1.085 0.276 ;
        RECT 1.499 0.252 1.541 0.294 ;
        RECT 1.803 0.252 1.845 0.294 ;
        RECT 0.587 0.325 0.629 0.367 ;
        RECT 0.891 0.326 0.933 0.368 ;
        RECT 1.043 0.326 1.085 0.368 ;
        RECT 1.499 0.344 1.541 0.386 ;
        RECT 1.499 0.436 1.541 0.478 ;
      LAYER M1 ;
        RECT 1.495 0.03 1.545 0.498 ;
        RECT 0.887 0.03 0.937 0.388 ;
        RECT 1.039 0.03 1.089 0.388 ;
        RECT 0.583 0.03 0.633 0.387 ;
        RECT 1.799 0.03 1.849 0.329 ;
        RECT 0 -0.03 2.128 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.283 1.38 0.325 1.422 ;
      RECT 0.283 1.472 0.325 1.514 ;
      RECT 1.347 0.251 1.389 0.293 ;
      RECT 0.283 1.38 0.325 1.422 ;
      RECT 1.347 0.343 1.389 0.385 ;
      RECT 0.283 0.351 0.325 0.393 ;
      RECT 0.283 1.472 0.325 1.514 ;
      RECT 0.511 0.551 0.553 0.593 ;
      RECT 0.283 1.288 0.325 1.33 ;
      RECT 0.283 1.288 0.325 1.33 ;
      RECT 1.347 1.481 1.389 1.523 ;
      RECT 0.739 0.164 0.781 0.206 ;
      RECT 1.347 1.389 1.389 1.431 ;
      RECT 1.347 1.205 1.389 1.247 ;
      RECT 0.283 1.196 0.325 1.238 ;
      RECT 1.347 1.389 1.389 1.431 ;
      RECT 1.347 1.297 1.389 1.339 ;
      RECT 1.347 1.297 1.389 1.339 ;
      RECT 1.727 0.614 1.769 0.656 ;
      RECT 1.575 0.614 1.617 0.656 ;
      RECT 0.739 1.06 0.781 1.102 ;
      RECT 0.283 1.104 0.325 1.146 ;
      RECT 0.739 0.348 0.781 0.39 ;
      RECT 0.739 0.256 0.781 0.298 ;
      RECT 0.283 0.167 0.325 0.209 ;
      RECT 1.347 1.481 1.389 1.523 ;
      RECT 0.283 0.259 0.325 0.301 ;
      RECT 1.347 0.159 1.389 0.201 ;
      RECT 1.119 0.968 1.161 1.01 ;
    LAYER M1 ;
      RECT 1.115 0.746 1.293 0.796 ;
      RECT 0.507 0.514 1.293 0.564 ;
      RECT 1.243 0.564 1.293 0.746 ;
      RECT 1.115 0.796 1.165 0.98 ;
      RECT 0.735 1.014 1.164 1.03 ;
      RECT 0.735 0.98 1.165 1.014 ;
      RECT 0.507 0.564 0.557 0.613 ;
      RECT 0.507 0.509 0.557 0.514 ;
      RECT 0.735 1.03 0.785 1.122 ;
      RECT 0.735 0.144 0.785 0.514 ;
      RECT 1.343 0.61 1.789 0.66 ;
      RECT 0.279 1.172 1.588 1.222 ;
      RECT 1.538 0.66 1.588 1.172 ;
      RECT 0.097 0.424 0.147 0.894 ;
      RECT 0.097 0.374 0.329 0.424 ;
      RECT 0.279 0.138 0.329 0.374 ;
      RECT 0.097 0.894 0.329 0.944 ;
      RECT 0.279 1.222 0.329 1.549 ;
      RECT 0.279 0.944 0.329 1.172 ;
      RECT 1.343 1.222 1.393 1.55 ;
      RECT 1.343 0.124 1.393 0.61 ;
    LAYER PO ;
      RECT 1.125 0.072 1.155 0.711 ;
      RECT 1.885 0.058 1.915 1.596 ;
      RECT 1.733 0.072 1.763 1.604 ;
      RECT 1.581 0.072 1.611 1.61 ;
      RECT 0.517 0.933 0.547 1.609 ;
      RECT 1.429 0.072 1.459 1.61 ;
      RECT 1.277 0.072 1.307 1.61 ;
      RECT 0.973 0.072 1.003 1.61 ;
      RECT 1.125 0.934 1.155 1.61 ;
      RECT 0.821 0.072 0.851 1.61 ;
      RECT 0.517 0.071 0.547 0.627 ;
      RECT 0.669 0.071 0.699 1.609 ;
      RECT 0.213 0.071 0.243 1.609 ;
      RECT 0.365 0.069 0.395 1.609 ;
      RECT 2.037 0.058 2.067 1.596 ;
      RECT 0.061 0.071 0.091 1.609 ;
    LAYER NWELL ;
      RECT -0.115 0.679 2.243 1.773 ;
  END
END MUX21X2_RVT

MACRO OA22X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.271 0.81 0.421 0.817 ;
        RECT 0.249 0.71 0.421 0.81 ;
        RECT 0.249 0.701 0.359 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0216 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.482 0.553 1.524 ;
      LAYER M1 ;
        RECT 0.401 1.571 0.511 1.577 ;
        RECT 0.401 1.461 0.573 1.571 ;
        RECT 0.426 1.46 0.573 1.461 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0216 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.744 0.857 0.786 ;
      LAYER M1 ;
        RECT 0.811 1.002 0.968 1.139 ;
        RECT 0.811 0.715 0.861 1.002 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0216 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.747 0.705 0.789 ;
      LAYER M1 ;
        RECT 0.56 0.963 0.709 0.986 ;
        RECT 0.553 0.854 0.709 0.963 ;
        RECT 0.659 0.723 0.709 0.854 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0216 ;
  END A4
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.043 0.239 1.085 0.281 ;
        RECT 1.347 0.239 1.389 0.281 ;
        RECT 1.043 0.331 1.085 0.373 ;
        RECT 1.347 0.331 1.389 0.373 ;
        RECT 1.043 0.423 1.085 0.465 ;
        RECT 1.347 0.423 1.389 0.465 ;
        RECT 1.347 0.987 1.389 1.029 ;
        RECT 1.347 1.079 1.389 1.121 ;
        RECT 1.347 1.171 1.389 1.213 ;
        RECT 1.347 1.263 1.389 1.305 ;
        RECT 1.347 1.355 1.389 1.397 ;
        RECT 1.043 1.395 1.085 1.437 ;
        RECT 1.043 1.487 1.085 1.529 ;
      LAYER M1 ;
        RECT 1.039 1.389 1.089 1.558 ;
        RECT 1.343 1.389 1.393 1.426 ;
        RECT 1.039 1.339 1.393 1.389 ;
        RECT 1.343 1.006 1.393 1.339 ;
        RECT 1.343 0.956 1.532 1.006 ;
        RECT 1.482 0.542 1.532 0.956 ;
        RECT 1.039 0.53 1.532 0.542 ;
        RECT 1.039 0.492 1.607 0.53 ;
        RECT 1.039 0.188 1.089 0.492 ;
        RECT 1.343 0.188 1.393 0.492 ;
        RECT 1.447 0.392 1.607 0.492 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.079 0.325 1.121 ;
        RECT 0.283 1.171 0.325 1.213 ;
        RECT 0.283 1.263 0.325 1.305 ;
        RECT 0.283 1.355 0.325 1.397 ;
        RECT 0.891 1.355 0.933 1.397 ;
        RECT 1.195 1.489 1.237 1.531 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.672 1.702 ;
        RECT 0.279 0.958 0.329 1.642 ;
        RECT 0.887 1.335 0.937 1.642 ;
        RECT 1.191 1.461 1.241 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.195 0.203 1.237 0.245 ;
        RECT 0.435 0.239 0.477 0.281 ;
        RECT 1.195 0.295 1.237 0.337 ;
        RECT 0.435 0.331 0.477 0.373 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.512 ;
        RECT 1.191 0.03 1.241 0.399 ;
        RECT 0 -0.03 1.672 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.231 0.681 1.317 0.699 ;
      RECT 1.231 0.613 1.317 0.631 ;
      RECT 0.735 0.631 1.317 0.663 ;
      RECT 1.07 0.663 1.317 0.681 ;
      RECT 1.07 0.681 1.156 0.699 ;
      RECT 1.079 0.699 1.129 1.226 ;
      RECT 0.583 1.226 1.129 1.276 ;
      RECT 0.735 0.613 1.156 0.631 ;
      RECT 0.735 0.212 0.785 0.613 ;
      RECT 0.583 1.276 0.633 1.393 ;
      RECT 0.583 1.106 0.633 1.226 ;
      RECT 0.583 0.095 0.937 0.145 ;
      RECT 0.887 0.145 0.937 0.504 ;
      RECT 0.583 0.145 0.633 0.598 ;
      RECT 0.279 0.598 0.633 0.648 ;
      RECT 0.279 0.178 0.329 0.598 ;
    LAYER PO ;
      RECT 1.429 0.101 1.459 1.469 ;
      RECT 0.821 0.101 0.851 1.469 ;
      RECT 0.669 0.101 0.699 1.469 ;
      RECT 1.125 0.069 1.155 1.608 ;
      RECT 0.365 0.101 0.395 1.469 ;
      RECT 1.581 0.101 1.611 1.469 ;
      RECT 0.517 0.101 0.547 1.567 ;
      RECT 1.277 0.069 1.307 1.608 ;
      RECT 0.973 0.101 1.003 1.469 ;
      RECT 0.061 0.101 0.091 1.469 ;
      RECT 0.213 0.101 0.243 1.469 ;
    LAYER CO ;
      RECT 1.271 0.635 1.313 0.677 ;
      RECT 0.587 1.322 0.629 1.364 ;
      RECT 0.587 1.23 0.629 1.272 ;
      RECT 0.587 1.138 0.629 1.18 ;
      RECT 1.119 0.635 1.161 0.677 ;
      RECT 0.587 0.239 0.629 0.281 ;
      RECT 0.587 0.331 0.629 0.373 ;
      RECT 0.283 0.239 0.325 0.281 ;
      RECT 0.739 0.239 0.781 0.281 ;
      RECT 0.891 0.331 0.933 0.373 ;
      RECT 0.891 0.239 0.933 0.281 ;
      RECT 0.283 0.331 0.325 0.373 ;
      RECT 0.739 0.331 0.781 0.373 ;
    LAYER NWELL ;
      RECT -0.135 0.679 1.788 1.787 ;
  END
END OA22X2_RVT

MACRO OAI21X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.271 0.81 0.421 0.817 ;
        RECT 0.249 0.717 0.421 0.81 ;
        RECT 0.249 0.701 0.359 0.717 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.482 0.553 1.524 ;
      LAYER M1 ;
        RECT 0.401 1.571 0.511 1.576 ;
        RECT 0.401 1.465 0.573 1.571 ;
        RECT 0.426 1.46 0.573 1.465 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.827 0.857 0.869 ;
      LAYER M1 ;
        RECT 0.712 0.962 0.861 0.986 ;
        RECT 0.705 0.853 0.861 0.962 ;
        RECT 0.811 0.807 0.861 0.853 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0138 ;
  END A3
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.499 0.239 1.541 0.281 ;
        RECT 1.499 0.331 1.541 0.373 ;
        RECT 1.499 0.423 1.541 0.465 ;
        RECT 1.499 0.987 1.541 1.029 ;
        RECT 1.499 1.079 1.541 1.121 ;
        RECT 1.499 1.171 1.541 1.213 ;
        RECT 1.499 1.263 1.541 1.305 ;
        RECT 1.499 1.355 1.541 1.397 ;
      LAYER M1 ;
        RECT 1.495 1.006 1.545 1.426 ;
        RECT 1.495 0.956 1.684 1.006 ;
        RECT 1.634 0.542 1.684 0.956 ;
        RECT 1.495 0.53 1.684 0.542 ;
        RECT 1.495 0.492 1.743 0.53 ;
        RECT 1.495 0.188 1.545 0.492 ;
        RECT 1.607 0.392 1.743 0.492 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 0.987 0.325 1.029 ;
        RECT 0.283 1.079 0.325 1.121 ;
        RECT 0.283 1.171 0.325 1.213 ;
        RECT 1.347 1.171 1.389 1.213 ;
        RECT 0.283 1.263 0.325 1.305 ;
        RECT 0.891 1.263 0.933 1.305 ;
        RECT 1.347 1.263 1.389 1.305 ;
        RECT 0.283 1.355 0.325 1.397 ;
        RECT 0.891 1.355 0.933 1.397 ;
        RECT 1.347 1.355 1.389 1.397 ;
        RECT 1.043 1.461 1.085 1.503 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.824 1.702 ;
        RECT 0.279 0.958 0.329 1.642 ;
        RECT 0.887 1.243 0.937 1.642 ;
        RECT 1.039 1.414 1.089 1.642 ;
        RECT 1.343 1.133 1.393 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.043 0.146 1.085 0.188 ;
        RECT 1.347 0.203 1.389 0.245 ;
        RECT 0.435 0.239 0.477 0.281 ;
        RECT 1.347 0.295 1.389 0.337 ;
        RECT 0.435 0.331 0.477 0.373 ;
        RECT 0.435 0.423 0.477 0.465 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.512 ;
        RECT 1.343 0.03 1.393 0.399 ;
        RECT 1.039 0.03 1.089 0.234 ;
        RECT 0 -0.03 1.824 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.079 0.785 1.165 0.803 ;
      RECT 1.079 0.717 1.165 0.735 ;
      RECT 0.913 0.755 1.165 0.785 ;
      RECT 0.887 0.735 1.165 0.755 ;
      RECT 0.887 0.705 0.963 0.735 ;
      RECT 0.583 1.13 0.963 1.18 ;
      RECT 0.887 0.181 0.937 0.705 ;
      RECT 0.913 0.785 0.963 1.13 ;
      RECT 0.583 1.18 0.633 1.393 ;
      RECT 0.583 1.106 0.633 1.13 ;
      RECT 0.735 1.18 0.785 1.393 ;
      RECT 0.735 1.106 0.785 1.13 ;
      RECT 1.231 0.631 1.48 0.681 ;
      RECT 1.383 0.681 1.469 0.699 ;
      RECT 1.383 0.613 1.469 0.631 ;
      RECT 1.231 0.681 1.281 0.956 ;
      RECT 1.231 0.542 1.281 0.631 ;
      RECT 1.191 0.492 1.281 0.542 ;
      RECT 1.191 0.089 1.241 0.492 ;
      RECT 1.191 0.956 1.281 1.006 ;
      RECT 1.191 1.006 1.241 1.555 ;
      RECT 0.279 0.598 0.633 0.648 ;
      RECT 0.735 0.181 0.785 0.412 ;
      RECT 0.583 0.412 0.785 0.462 ;
      RECT 0.583 0.462 0.633 0.598 ;
      RECT 0.583 0.181 0.633 0.412 ;
      RECT 0.279 0.178 0.329 0.598 ;
    LAYER PO ;
      RECT 0.973 0.101 1.003 1.469 ;
      RECT 1.125 0.054 1.155 1.608 ;
      RECT 0.365 0.101 0.395 1.469 ;
      RECT 0.821 0.101 0.851 1.469 ;
      RECT 1.581 0.101 1.611 1.469 ;
      RECT 1.733 0.101 1.763 1.469 ;
      RECT 0.061 0.101 0.091 1.469 ;
      RECT 1.277 0.101 1.307 1.469 ;
      RECT 1.429 0.069 1.459 1.608 ;
      RECT 0.517 0.101 0.547 1.567 ;
      RECT 0.213 0.101 0.243 1.469 ;
      RECT 0.669 0.101 0.699 1.469 ;
    LAYER CO ;
      RECT 0.587 0.331 0.629 0.373 ;
      RECT 1.423 0.635 1.465 0.677 ;
      RECT 0.891 0.211 0.933 0.253 ;
      RECT 0.891 0.303 0.933 0.345 ;
      RECT 0.283 0.239 0.325 0.281 ;
      RECT 1.119 0.739 1.161 0.781 ;
      RECT 0.739 1.23 0.781 1.272 ;
      RECT 0.739 1.322 0.781 1.364 ;
      RECT 1.195 1.454 1.237 1.496 ;
      RECT 0.587 0.423 0.629 0.465 ;
      RECT 0.283 0.423 0.325 0.465 ;
      RECT 0.283 0.331 0.325 0.373 ;
      RECT 0.739 0.303 0.781 0.345 ;
      RECT 0.739 0.211 0.781 0.253 ;
      RECT 0.587 1.23 0.629 1.272 ;
      RECT 0.587 1.322 0.629 1.364 ;
      RECT 0.587 1.138 0.629 1.18 ;
      RECT 1.195 0.145 1.237 0.187 ;
      RECT 0.587 0.239 0.629 0.281 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.939 1.787 ;
  END
END OAI21X1_RVT

MACRO AO21X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.897 0.553 0.939 ;
      LAYER M1 ;
        RECT 0.491 0.857 0.663 0.967 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0243 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.732 0.401 0.774 ;
      LAYER M1 ;
        RECT 0.249 0.705 0.421 0.815 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0243 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.124 0.857 0.166 ;
      LAYER M1 ;
        RECT 0.705 0.097 0.877 0.207 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0225 ;
  END A3
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.043 0.18 1.085 0.222 ;
        RECT 1.347 0.18 1.389 0.222 ;
        RECT 1.043 0.272 1.085 0.314 ;
        RECT 1.347 0.272 1.389 0.314 ;
        RECT 1.043 0.364 1.085 0.406 ;
        RECT 1.347 0.364 1.389 0.406 ;
        RECT 1.043 0.456 1.085 0.498 ;
        RECT 1.347 0.456 1.389 0.498 ;
        RECT 1.043 0.764 1.085 0.806 ;
        RECT 1.347 0.838 1.389 0.88 ;
        RECT 1.043 0.856 1.085 0.898 ;
        RECT 1.347 0.93 1.389 0.972 ;
        RECT 1.043 0.948 1.085 0.99 ;
        RECT 1.347 1.022 1.389 1.064 ;
        RECT 1.043 1.04 1.085 1.082 ;
        RECT 1.347 1.114 1.389 1.156 ;
        RECT 1.347 1.206 1.389 1.248 ;
        RECT 1.347 1.298 1.389 1.34 ;
        RECT 1.347 1.39 1.389 1.432 ;
        RECT 1.347 1.482 1.389 1.524 ;
      LAYER M1 ;
        RECT 1.344 1.119 1.394 1.544 ;
        RECT 1.313 1.009 1.423 1.119 ;
        RECT 1.039 0.794 1.089 1.102 ;
        RECT 1.344 0.75 1.394 1.009 ;
        RECT 1.01 0.744 1.089 0.794 ;
        RECT 1.344 0.7 1.432 0.75 ;
        RECT 1.01 0.518 1.06 0.744 ;
        RECT 1.382 0.518 1.432 0.7 ;
        RECT 1.01 0.468 1.432 0.518 ;
        RECT 1.039 0.16 1.089 0.468 ;
        RECT 1.344 0.16 1.394 0.468 ;
    END
    ANTENNADIFFAREA 0.2484 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.14 0.325 1.182 ;
        RECT 0.283 1.232 0.325 1.274 ;
        RECT 0.587 1.232 0.629 1.274 ;
        RECT 1.195 1.308 1.237 1.35 ;
        RECT 0.283 1.324 0.325 1.366 ;
        RECT 0.587 1.324 0.629 1.366 ;
        RECT 1.195 1.4 1.237 1.442 ;
        RECT 0.283 1.416 0.325 1.458 ;
        RECT 0.587 1.416 0.629 1.458 ;
        RECT 1.195 1.492 1.237 1.534 ;
        RECT 0.283 1.508 0.325 1.55 ;
        RECT 0.587 1.508 0.629 1.55 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.672 1.702 ;
        RECT 0.279 1.12 0.329 1.642 ;
        RECT 0.583 1.212 0.633 1.642 ;
        RECT 1.191 1.288 1.241 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.195 0.134 1.237 0.176 ;
        RECT 1.195 0.226 1.237 0.268 ;
        RECT 1.195 0.318 1.237 0.36 ;
        RECT 0.283 0.415 0.325 0.457 ;
        RECT 0.739 0.415 0.781 0.457 ;
        RECT 0.283 0.507 0.325 0.549 ;
        RECT 0.739 0.507 0.781 0.549 ;
      LAYER M1 ;
        RECT 0.279 0.345 0.329 0.569 ;
        RECT 0.735 0.345 0.785 0.569 ;
        RECT 0.279 0.295 0.785 0.345 ;
        RECT 1.191 0.03 1.241 0.38 ;
        RECT 0.279 0.03 0.329 0.295 ;
        RECT 0 -0.03 1.672 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.115 0.568 1.317 0.65 ;
      RECT 1.198 0.65 1.248 1.152 ;
      RECT 0.887 1.152 1.248 1.202 ;
      RECT 0.887 1.202 0.937 1.575 ;
      RECT 0.583 0.651 0.937 0.701 ;
      RECT 0.887 0.701 0.937 1.152 ;
      RECT 0.887 0.395 0.937 0.651 ;
      RECT 0.583 0.395 0.633 0.651 ;
      RECT 0.735 1.127 0.785 1.57 ;
      RECT 0.431 1.077 0.785 1.127 ;
      RECT 0.431 1.127 0.481 1.575 ;
    LAYER PO ;
      RECT 1.429 0.056 1.459 1.597 ;
      RECT 0.517 0.071 0.547 1.62 ;
      RECT 1.581 0.056 1.611 1.597 ;
      RECT 0.061 0.064 0.091 1.613 ;
      RECT 0.669 0.071 0.699 1.62 ;
      RECT 0.365 0.066 0.395 1.62 ;
      RECT 0.821 0.066 0.851 1.62 ;
      RECT 1.277 0.052 1.307 1.604 ;
      RECT 0.973 0.064 1.003 1.613 ;
      RECT 1.125 0.064 1.155 1.604 ;
      RECT 0.213 0.064 0.243 1.613 ;
    LAYER CO ;
      RECT 0.435 1.508 0.477 1.55 ;
      RECT 0.891 0.507 0.933 0.549 ;
      RECT 0.891 1.508 0.933 1.55 ;
      RECT 1.271 0.588 1.313 0.63 ;
      RECT 0.435 1.14 0.477 1.182 ;
      RECT 0.739 1.14 0.781 1.182 ;
      RECT 0.739 1.232 0.781 1.274 ;
      RECT 0.891 1.14 0.933 1.182 ;
      RECT 0.891 1.232 0.933 1.274 ;
      RECT 0.891 0.415 0.933 0.457 ;
      RECT 0.891 1.416 0.933 1.458 ;
      RECT 0.891 1.324 0.933 1.366 ;
      RECT 0.891 1.048 0.933 1.09 ;
      RECT 0.739 1.416 0.781 1.458 ;
      RECT 0.587 0.507 0.629 0.549 ;
      RECT 0.587 0.415 0.629 0.457 ;
      RECT 0.435 1.232 0.477 1.274 ;
      RECT 0.739 1.508 0.781 1.55 ;
      RECT 1.119 0.588 1.161 0.63 ;
      RECT 0.739 1.324 0.781 1.366 ;
      RECT 0.435 1.324 0.477 1.366 ;
      RECT 0.435 1.416 0.477 1.458 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.787 1.773 ;
  END
END AO21X2_RVT

MACRO OA222X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.128 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.271 0.81 0.421 0.817 ;
        RECT 0.249 0.71 0.421 0.81 ;
        RECT 0.249 0.701 0.359 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.482 0.553 1.524 ;
      LAYER M1 ;
        RECT 0.401 1.571 0.511 1.577 ;
        RECT 0.401 1.461 0.573 1.571 ;
        RECT 0.426 1.46 0.573 1.461 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.807 0.857 0.849 ;
      LAYER M1 ;
        RECT 0.811 1.002 0.968 1.139 ;
        RECT 0.811 0.772 0.861 1.002 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.739 0.705 0.781 ;
      LAYER M1 ;
        RECT 0.56 0.963 0.709 0.986 ;
        RECT 0.553 0.854 0.709 0.963 ;
        RECT 0.659 0.713 0.709 0.854 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.119 0.739 1.161 0.781 ;
      LAYER M1 ;
        RECT 1.115 0.675 1.165 0.808 ;
        RECT 1.023 0.658 1.165 0.675 ;
        RECT 1.009 0.601 1.165 0.658 ;
        RECT 1.009 0.549 1.123 0.601 ;
        RECT 1.023 0.541 1.123 0.549 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A5
  PIN A6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.271 1.49 1.313 1.532 ;
      LAYER M1 ;
        RECT 1.171 1.485 1.339 1.535 ;
        RECT 1.171 1.281 1.221 1.485 ;
        RECT 1.171 1.266 1.28 1.281 ;
        RECT 1.16 1.157 1.28 1.266 ;
        RECT 1.171 1.146 1.28 1.157 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A6
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.499 0.239 1.541 0.281 ;
        RECT 1.803 0.239 1.845 0.281 ;
        RECT 1.499 0.331 1.541 0.373 ;
        RECT 1.803 0.331 1.845 0.373 ;
        RECT 1.499 0.423 1.541 0.465 ;
        RECT 1.803 0.423 1.845 0.465 ;
        RECT 1.499 0.987 1.541 1.029 ;
        RECT 1.803 0.987 1.845 1.029 ;
        RECT 1.499 1.079 1.541 1.121 ;
        RECT 1.803 1.079 1.845 1.121 ;
        RECT 1.499 1.171 1.541 1.213 ;
        RECT 1.803 1.171 1.845 1.213 ;
        RECT 1.499 1.263 1.541 1.305 ;
        RECT 1.803 1.263 1.845 1.305 ;
        RECT 1.499 1.355 1.541 1.397 ;
        RECT 1.803 1.355 1.845 1.397 ;
      LAYER M1 ;
        RECT 1.495 1.006 1.545 1.426 ;
        RECT 1.799 1.006 1.849 1.426 ;
        RECT 1.495 0.956 1.988 1.006 ;
        RECT 1.938 0.542 1.988 0.956 ;
        RECT 1.495 0.53 1.988 0.542 ;
        RECT 1.495 0.492 2.063 0.53 ;
        RECT 1.495 0.188 1.545 0.492 ;
        RECT 1.799 0.188 1.849 0.492 ;
        RECT 1.903 0.392 2.063 0.492 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.079 0.325 1.121 ;
        RECT 0.283 1.171 0.325 1.213 ;
        RECT 1.651 1.171 1.693 1.213 ;
        RECT 0.283 1.263 0.325 1.305 ;
        RECT 1.651 1.263 1.693 1.305 ;
        RECT 0.283 1.355 0.325 1.397 ;
        RECT 0.891 1.355 0.933 1.397 ;
        RECT 1.043 1.355 1.085 1.397 ;
        RECT 1.651 1.355 1.693 1.397 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 2.128 1.702 ;
        RECT 0.279 0.958 0.329 1.642 ;
        RECT 0.887 1.335 0.937 1.642 ;
        RECT 1.039 1.333 1.089 1.642 ;
        RECT 1.647 1.133 1.697 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 1.651 0.203 1.693 0.245 ;
        RECT 0.435 0.239 0.477 0.281 ;
        RECT 1.651 0.295 1.693 0.337 ;
        RECT 0.435 0.331 0.477 0.373 ;
        RECT 0.435 0.423 0.477 0.465 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.512 ;
        RECT 1.647 0.03 1.697 0.399 ;
        RECT 0 -0.03 2.128 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.687 0.681 1.773 0.699 ;
      RECT 1.687 0.613 1.773 0.631 ;
      RECT 1.343 0.631 1.773 0.681 ;
      RECT 0.583 1.263 0.633 1.393 ;
      RECT 0.583 1.106 0.633 1.213 ;
      RECT 1.526 0.681 1.612 0.699 ;
      RECT 1.526 0.613 1.612 0.631 ;
      RECT 1.039 0.903 1.393 0.953 ;
      RECT 1.191 0.483 1.393 0.533 ;
      RECT 1.343 0.953 1.393 1.38 ;
      RECT 1.191 0.211 1.241 0.483 ;
      RECT 1.343 0.681 1.393 0.903 ;
      RECT 1.343 0.533 1.393 0.631 ;
      RECT 1.039 0.953 1.089 1.213 ;
      RECT 0.583 1.213 1.089 1.263 ;
      RECT 1.039 0.148 1.089 0.431 ;
      RECT 0.735 0.098 1.393 0.148 ;
      RECT 1.343 0.148 1.393 0.432 ;
      RECT 0.735 0.148 0.785 0.501 ;
      RECT 0.279 0.598 0.937 0.648 ;
      RECT 0.583 0.181 0.633 0.598 ;
      RECT 0.887 0.208 0.937 0.598 ;
      RECT 0.279 0.178 0.329 0.598 ;
    LAYER PO ;
      RECT 1.581 0.069 1.611 1.608 ;
      RECT 1.733 0.069 1.763 1.608 ;
      RECT 0.821 0.101 0.851 1.469 ;
      RECT 0.669 0.101 0.699 1.469 ;
      RECT 0.517 0.101 0.547 1.567 ;
      RECT 0.213 0.101 0.243 1.469 ;
      RECT 1.277 0.101 1.307 1.567 ;
      RECT 1.125 0.101 1.155 1.469 ;
      RECT 0.365 0.101 0.395 1.469 ;
      RECT 1.429 0.101 1.459 1.469 ;
      RECT 1.885 0.101 1.915 1.469 ;
      RECT 2.037 0.101 2.067 1.469 ;
      RECT 0.061 0.101 0.091 1.469 ;
      RECT 0.973 0.101 1.003 1.469 ;
    LAYER CO ;
      RECT 0.587 1.138 0.629 1.18 ;
      RECT 1.575 0.635 1.617 0.677 ;
      RECT 0.587 1.322 0.629 1.364 ;
      RECT 0.587 1.23 0.629 1.272 ;
      RECT 1.347 1.289 1.389 1.331 ;
      RECT 1.347 1.197 1.389 1.239 ;
      RECT 1.043 0.27 1.085 0.312 ;
      RECT 1.043 0.362 1.085 0.404 ;
      RECT 0.891 0.239 0.933 0.281 ;
      RECT 0.891 0.331 0.933 0.373 ;
      RECT 1.043 0.178 1.085 0.22 ;
      RECT 0.739 0.331 0.781 0.373 ;
      RECT 0.587 0.239 0.629 0.281 ;
      RECT 0.283 0.239 0.325 0.281 ;
      RECT 0.739 0.423 0.781 0.465 ;
      RECT 0.739 0.239 0.781 0.281 ;
      RECT 1.195 0.362 1.237 0.404 ;
      RECT 0.587 0.423 0.629 0.465 ;
      RECT 1.347 0.27 1.389 0.312 ;
      RECT 1.347 0.362 1.389 0.404 ;
      RECT 1.347 0.178 1.389 0.22 ;
      RECT 1.727 0.635 1.769 0.677 ;
      RECT 0.283 0.423 0.325 0.465 ;
      RECT 0.283 0.331 0.325 0.373 ;
      RECT 1.195 0.27 1.237 0.312 ;
      RECT 0.891 0.423 0.933 0.465 ;
      RECT 0.587 0.331 0.629 0.373 ;
    LAYER NWELL ;
      RECT -0.135 0.679 2.244 1.787 ;
  END
END OA222X2_RVT

MACRO OR2X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.368 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.664 0.401 0.706 ;
      LAYER M1 ;
        RECT 0.249 0.857 0.405 0.967 ;
        RECT 0.355 0.644 0.405 0.857 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0306 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.664 0.553 0.706 ;
      LAYER M1 ;
        RECT 0.505 0.642 0.663 0.815 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0306 ;
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.891 0.228 0.933 0.27 ;
        RECT 0.891 0.32 0.933 0.362 ;
        RECT 0.891 0.412 0.933 0.454 ;
        RECT 0.891 0.506 0.933 0.548 ;
        RECT 0.891 0.817 0.933 0.859 ;
        RECT 0.891 0.909 0.933 0.951 ;
        RECT 0.891 1.001 0.933 1.043 ;
        RECT 0.891 1.093 0.933 1.135 ;
        RECT 0.891 1.185 0.933 1.227 ;
        RECT 0.891 1.277 0.933 1.319 ;
        RECT 0.891 1.371 0.933 1.413 ;
        RECT 0.891 1.463 0.933 1.505 ;
      LAYER M1 ;
        RECT 0.887 0.89 0.937 1.525 ;
        RECT 0.887 0.84 1.157 0.89 ;
        RECT 0.887 0.797 0.937 0.84 ;
        RECT 1.107 0.663 1.157 0.84 ;
        RECT 1.107 0.595 1.271 0.663 ;
        RECT 0.887 0.545 1.271 0.595 ;
        RECT 0.887 0.208 0.937 0.545 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.043 1.016 1.085 1.058 ;
        RECT 0.283 1.107 0.325 1.149 ;
        RECT 0.739 1.107 0.781 1.149 ;
        RECT 1.043 1.108 1.085 1.15 ;
        RECT 0.283 1.2 0.325 1.242 ;
        RECT 0.739 1.2 0.781 1.242 ;
        RECT 1.043 1.2 1.085 1.242 ;
        RECT 0.283 1.292 0.325 1.334 ;
        RECT 0.739 1.292 0.781 1.334 ;
        RECT 1.043 1.292 1.085 1.334 ;
        RECT 0.283 1.386 0.325 1.428 ;
        RECT 0.739 1.386 0.781 1.428 ;
        RECT 1.043 1.386 1.085 1.428 ;
        RECT 0.283 1.478 0.325 1.52 ;
        RECT 0.739 1.478 0.781 1.52 ;
        RECT 1.043 1.478 1.085 1.52 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.368 1.702 ;
        RECT 0.279 1.087 0.329 1.642 ;
        RECT 0.735 1.087 0.785 1.642 ;
        RECT 1.039 0.996 1.089 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 0.739 0.228 0.781 0.27 ;
        RECT 1.043 0.228 1.085 0.27 ;
        RECT 0.739 0.32 0.781 0.362 ;
        RECT 1.043 0.32 1.085 0.362 ;
        RECT 0.435 0.337 0.477 0.379 ;
        RECT 1.043 0.412 1.085 0.454 ;
      LAYER M1 ;
        RECT 1.039 0.03 1.089 0.474 ;
        RECT 0.431 0.03 0.481 0.399 ;
        RECT 0.735 0.03 0.785 0.382 ;
        RECT 0 -0.03 1.368 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.781 0.66 1.029 0.71 ;
      RECT 0.583 0.933 0.806 0.983 ;
      RECT 0.756 0.511 0.806 0.961 ;
      RECT 0.278 0.486 0.806 0.536 ;
      RECT 0.279 0.319 0.329 0.534 ;
      RECT 0.583 0.933 0.633 1.525 ;
      RECT 0.583 0.321 0.633 0.534 ;
    LAYER PO ;
      RECT 1.125 0.093 1.155 1.606 ;
      RECT 0.973 0.093 1.003 1.606 ;
      RECT 0.821 0.093 0.851 1.606 ;
      RECT 1.277 0.093 1.307 1.606 ;
      RECT 0.061 0.093 0.091 1.606 ;
      RECT 0.213 0.093 0.243 1.606 ;
      RECT 0.669 0.093 0.699 1.606 ;
      RECT 0.365 0.093 0.395 1.606 ;
      RECT 0.517 0.093 0.547 1.606 ;
    LAYER CO ;
      RECT 0.815 0.664 0.857 0.706 ;
      RECT 0.967 0.664 1.009 0.706 ;
      RECT 0.283 0.431 0.325 0.473 ;
      RECT 0.283 0.339 0.325 0.381 ;
      RECT 0.587 1.463 0.629 1.505 ;
      RECT 0.587 1.371 0.629 1.413 ;
      RECT 0.587 1.277 0.629 1.319 ;
      RECT 0.587 1.185 0.629 1.227 ;
      RECT 0.587 0.341 0.629 0.383 ;
      RECT 0.587 1.093 0.629 1.135 ;
      RECT 0.587 0.433 0.629 0.475 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.483 1.773 ;
  END
END OR2X2_RVT

MACRO AO221X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.808 0.401 0.85 ;
      LAYER M1 ;
        RECT 0.249 0.857 0.405 0.967 ;
        RECT 0.355 0.788 0.405 0.857 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.502 0.553 0.544 ;
      LAYER M1 ;
        RECT 0.401 0.498 0.573 0.548 ;
        RECT 0.401 0.359 0.451 0.498 ;
        RECT 0.401 0.249 0.511 0.359 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.112 0.857 0.154 ;
      LAYER M1 ;
        RECT 0.705 0.097 0.88 0.207 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.805 0.705 0.847 ;
      LAYER M1 ;
        RECT 0.553 1.009 0.663 1.119 ;
        RECT 0.606 0.851 0.656 1.009 ;
        RECT 0.606 0.801 0.725 0.851 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.119 0.777 1.161 0.819 ;
      LAYER M1 ;
        RECT 1.009 0.773 1.181 0.823 ;
        RECT 1.009 0.705 1.119 0.773 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END A5
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.347 0.194 1.389 0.236 ;
        RECT 1.651 0.194 1.693 0.236 ;
        RECT 1.347 0.286 1.389 0.328 ;
        RECT 1.651 0.286 1.693 0.328 ;
        RECT 1.347 0.378 1.389 0.42 ;
        RECT 1.651 0.378 1.693 0.42 ;
        RECT 1.347 0.47 1.389 0.512 ;
        RECT 1.651 0.47 1.693 0.512 ;
        RECT 1.347 0.778 1.389 0.82 ;
        RECT 1.651 0.778 1.693 0.82 ;
        RECT 1.347 0.87 1.389 0.912 ;
        RECT 1.651 0.87 1.693 0.912 ;
        RECT 1.347 0.962 1.389 1.004 ;
        RECT 1.651 0.962 1.693 1.004 ;
        RECT 1.347 1.054 1.389 1.096 ;
        RECT 1.651 1.054 1.693 1.096 ;
        RECT 1.651 1.146 1.693 1.188 ;
        RECT 1.651 1.238 1.693 1.28 ;
        RECT 1.651 1.33 1.693 1.372 ;
        RECT 1.651 1.422 1.693 1.464 ;
      LAYER M1 ;
        RECT 1.648 1.119 1.698 1.484 ;
        RECT 1.617 1.009 1.727 1.119 ;
        RECT 1.343 0.806 1.393 1.116 ;
        RECT 1.648 0.783 1.698 1.009 ;
        RECT 1.315 0.758 1.393 0.806 ;
        RECT 1.648 0.733 1.736 0.783 ;
        RECT 1.315 0.553 1.365 0.758 ;
        RECT 1.686 0.553 1.736 0.733 ;
        RECT 1.315 0.503 1.736 0.553 ;
        RECT 1.343 0.174 1.393 0.503 ;
        RECT 1.648 0.482 1.736 0.503 ;
        RECT 1.648 0.174 1.698 0.482 ;
    END
    ANTENNADIFFAREA 0.2484 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.499 1.312 1.541 1.354 ;
        RECT 1.499 1.404 1.541 1.446 ;
        RECT 0.435 1.407 0.477 1.449 ;
        RECT 1.499 1.496 1.541 1.538 ;
        RECT 0.435 1.499 0.477 1.541 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.976 1.702 ;
        RECT 0.431 1.387 0.481 1.642 ;
        RECT 1.495 1.284 1.545 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 1.499 0.148 1.541 0.19 ;
        RECT 0.587 0.212 0.629 0.254 ;
        RECT 1.499 0.24 1.541 0.282 ;
        RECT 0.587 0.304 0.629 0.346 ;
        RECT 1.499 0.332 1.541 0.374 ;
        RECT 1.043 0.335 1.085 0.377 ;
      LAYER M1 ;
        RECT 1.04 0.03 1.09 0.397 ;
        RECT 1.495 0.03 1.545 0.394 ;
        RECT 0.583 0.03 0.633 0.366 ;
        RECT 0 -0.03 1.976 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.419 0.603 1.621 0.685 ;
      RECT 1.19 1.184 1.543 1.234 ;
      RECT 1.493 0.685 1.543 1.184 ;
      RECT 0.279 0.276 0.329 0.598 ;
      RECT 0.279 0.632 0.937 0.648 ;
      RECT 0.887 0.648 0.937 0.917 ;
      RECT 0.887 0.273 0.937 0.582 ;
      RECT 0.887 0.917 1.24 0.967 ;
      RECT 1.19 1.234 1.24 1.571 ;
      RECT 1.19 0.967 1.24 1.184 ;
      RECT 1.192 0.309 1.242 0.582 ;
      RECT 0.279 0.598 1.242 0.632 ;
      RECT 0.887 0.582 1.242 0.598 ;
      RECT 0.735 1.021 1.089 1.071 ;
      RECT 1.039 1.071 1.089 1.571 ;
      RECT 0.735 1.071 0.785 1.237 ;
      RECT 0.583 1.337 0.633 1.564 ;
      RECT 0.279 1.287 0.937 1.337 ;
      RECT 0.887 1.337 0.937 1.571 ;
      RECT 0.279 1.337 0.329 1.571 ;
    LAYER PO ;
      RECT 1.733 0.07 1.763 1.611 ;
      RECT 1.277 0.075 1.307 1.616 ;
      RECT 1.429 0.078 1.459 1.618 ;
      RECT 1.581 0.066 1.611 1.618 ;
      RECT 1.885 0.07 1.915 1.611 ;
      RECT 0.669 0.072 0.699 1.621 ;
      RECT 0.517 0.072 0.547 1.621 ;
      RECT 0.365 0.067 0.395 1.621 ;
      RECT 0.061 0.072 0.091 1.621 ;
      RECT 0.973 0.076 1.003 1.621 ;
      RECT 0.821 0.072 0.851 1.621 ;
      RECT 0.213 0.072 0.243 1.621 ;
      RECT 1.125 0.076 1.155 1.621 ;
    LAYER CO ;
      RECT 0.891 0.293 0.933 0.335 ;
      RECT 1.195 1.141 1.237 1.183 ;
      RECT 0.283 0.296 0.325 0.338 ;
      RECT 0.891 1.417 0.933 1.459 ;
      RECT 1.195 1.325 1.237 1.367 ;
      RECT 1.195 1.417 1.237 1.459 ;
      RECT 1.195 1.233 1.237 1.275 ;
      RECT 1.195 1.509 1.237 1.551 ;
      RECT 1.043 1.509 1.085 1.551 ;
      RECT 1.195 0.337 1.237 0.379 ;
      RECT 0.587 1.502 0.629 1.544 ;
      RECT 1.043 1.325 1.085 1.367 ;
      RECT 1.043 1.417 1.085 1.459 ;
      RECT 1.423 0.623 1.465 0.665 ;
      RECT 1.575 0.623 1.617 0.665 ;
      RECT 0.891 1.325 0.933 1.367 ;
      RECT 0.283 1.417 0.325 1.459 ;
      RECT 0.283 1.509 0.325 1.551 ;
      RECT 0.739 1.175 0.781 1.217 ;
      RECT 0.739 1.083 0.781 1.125 ;
      RECT 0.587 1.41 0.629 1.452 ;
      RECT 0.587 1.318 0.629 1.36 ;
      RECT 0.283 1.325 0.325 1.367 ;
      RECT 0.283 0.388 0.325 0.43 ;
      RECT 0.891 0.385 0.933 0.427 ;
      RECT 0.891 1.509 0.933 1.551 ;
      RECT 1.043 1.233 1.085 1.275 ;
      RECT 1.043 1.141 1.085 1.183 ;
    LAYER NWELL ;
      RECT -0.115 0.679 2.091 1.773 ;
  END
END AO221X2_RVT

MACRO AOI22X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.744 0.401 0.786 ;
      LAYER M1 ;
        RECT 0.249 0.705 0.404 0.815 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0225 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.744 0.553 0.786 ;
      LAYER M1 ;
        RECT 0.401 1.009 0.557 1.119 ;
        RECT 0.507 0.724 0.557 1.009 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0225 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.108 0.857 0.15 ;
      LAYER M1 ;
        RECT 0.705 0.097 0.9 0.207 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0225 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.6 0.705 0.642 ;
      LAYER M1 ;
        RECT 0.553 0.553 0.708 0.663 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0225 ;
  END A4
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.347 0.18 1.389 0.222 ;
        RECT 1.651 0.18 1.693 0.222 ;
        RECT 1.347 0.272 1.389 0.314 ;
        RECT 1.651 0.272 1.693 0.314 ;
        RECT 1.347 0.364 1.389 0.406 ;
        RECT 1.651 0.364 1.693 0.406 ;
        RECT 1.347 0.456 1.389 0.498 ;
        RECT 1.651 0.456 1.693 0.498 ;
        RECT 1.347 0.764 1.389 0.806 ;
        RECT 1.651 0.764 1.693 0.806 ;
        RECT 1.347 0.856 1.389 0.898 ;
        RECT 1.651 0.856 1.693 0.898 ;
        RECT 1.347 0.948 1.389 0.99 ;
        RECT 1.651 0.948 1.693 0.99 ;
        RECT 1.347 1.04 1.389 1.082 ;
        RECT 1.651 1.04 1.693 1.082 ;
        RECT 1.651 1.132 1.693 1.174 ;
        RECT 1.651 1.224 1.693 1.266 ;
        RECT 1.651 1.316 1.693 1.358 ;
        RECT 1.651 1.408 1.693 1.45 ;
      LAYER M1 ;
        RECT 1.648 1.119 1.698 1.47 ;
        RECT 1.617 1.009 1.727 1.119 ;
        RECT 1.343 0.794 1.393 1.102 ;
        RECT 1.648 0.75 1.698 1.009 ;
        RECT 1.319 0.744 1.393 0.794 ;
        RECT 1.648 0.7 1.736 0.75 ;
        RECT 1.319 0.518 1.369 0.744 ;
        RECT 1.686 0.518 1.736 0.7 ;
        RECT 1.319 0.468 1.736 0.518 ;
        RECT 1.343 0.16 1.393 0.468 ;
        RECT 1.648 0.16 1.698 0.468 ;
    END
    ANTENNADIFFAREA 0.2484 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.043 1.041 1.085 1.083 ;
        RECT 1.043 1.133 1.085 1.175 ;
        RECT 1.043 1.225 1.085 1.267 ;
        RECT 1.043 1.317 1.085 1.359 ;
        RECT 1.499 1.39 1.541 1.432 ;
        RECT 0.435 1.407 0.477 1.449 ;
        RECT 1.043 1.409 1.085 1.451 ;
        RECT 1.499 1.482 1.541 1.524 ;
        RECT 0.435 1.499 0.477 1.541 ;
        RECT 1.043 1.501 1.085 1.543 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.976 1.702 ;
        RECT 0.431 1.387 0.481 1.642 ;
        RECT 1.039 1.021 1.089 1.642 ;
        RECT 1.495 1.37 1.545 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 1.499 0.134 1.541 0.176 ;
        RECT 0.587 0.2 0.629 0.242 ;
        RECT 1.043 0.204 1.085 0.246 ;
        RECT 1.499 0.226 1.541 0.268 ;
        RECT 0.587 0.292 0.629 0.334 ;
        RECT 1.043 0.296 1.085 0.338 ;
        RECT 1.043 0.388 1.085 0.43 ;
      LAYER M1 ;
        RECT 1.039 0.03 1.089 0.45 ;
        RECT 0.583 0.03 0.633 0.354 ;
        RECT 1.495 0.03 1.545 0.288 ;
        RECT 0 -0.03 1.976 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.419 0.568 1.621 0.65 ;
      RECT 1.495 0.65 1.545 1.229 ;
      RECT 1.191 1.229 1.545 1.279 ;
      RECT 1.191 0.606 1.269 0.656 ;
      RECT 1.191 1.279 1.241 1.563 ;
      RECT 1.191 1.105 1.241 1.229 ;
      RECT 1.191 1.055 1.269 1.105 ;
      RECT 1.191 0.184 1.241 0.606 ;
      RECT 1.219 0.656 1.269 1.055 ;
      RECT 1.116 0.712 1.166 0.813 ;
      RECT 0.735 0.813 1.166 0.863 ;
      RECT 0.279 0.261 0.329 0.422 ;
      RECT 0.735 0.863 0.785 1.237 ;
      RECT 0.758 0.472 0.808 0.813 ;
      RECT 0.887 0.264 0.937 0.422 ;
      RECT 0.279 0.422 0.937 0.472 ;
      RECT 0.583 1.337 0.633 1.571 ;
      RECT 0.279 1.287 0.937 1.337 ;
      RECT 0.887 1.337 0.937 1.571 ;
      RECT 0.279 1.337 0.329 1.571 ;
    LAYER PO ;
      RECT 1.733 0.056 1.763 1.597 ;
      RECT 0.669 0.072 0.699 1.621 ;
      RECT 0.517 0.072 0.547 1.621 ;
      RECT 0.365 0.067 0.395 1.621 ;
      RECT 0.061 0.072 0.091 1.621 ;
      RECT 0.973 0.076 1.003 1.621 ;
      RECT 0.821 0.072 0.851 1.621 ;
      RECT 0.213 0.072 0.243 1.621 ;
      RECT 1.277 0.076 1.307 1.621 ;
      RECT 1.581 0.052 1.611 1.604 ;
      RECT 1.885 0.056 1.915 1.597 ;
      RECT 1.429 0.064 1.459 1.604 ;
      RECT 1.125 0.059 1.155 1.613 ;
    LAYER CO ;
      RECT 1.575 0.588 1.617 0.63 ;
      RECT 1.423 0.588 1.465 0.63 ;
      RECT 1.195 1.409 1.237 1.451 ;
      RECT 1.195 1.501 1.237 1.543 ;
      RECT 1.195 1.317 1.237 1.359 ;
      RECT 1.195 1.225 1.237 1.267 ;
      RECT 1.195 1.133 1.237 1.175 ;
      RECT 0.739 1.175 0.781 1.217 ;
      RECT 0.739 1.083 0.781 1.125 ;
      RECT 0.587 1.417 0.629 1.459 ;
      RECT 0.587 1.325 0.629 1.367 ;
      RECT 0.891 1.417 0.933 1.459 ;
      RECT 0.891 0.376 0.933 0.418 ;
      RECT 0.283 1.417 0.325 1.459 ;
      RECT 0.891 0.284 0.933 0.326 ;
      RECT 0.283 0.281 0.325 0.323 ;
      RECT 0.283 0.373 0.325 0.415 ;
      RECT 0.891 1.325 0.933 1.367 ;
      RECT 0.891 1.509 0.933 1.551 ;
      RECT 0.283 1.325 0.325 1.367 ;
      RECT 0.283 1.509 0.325 1.551 ;
      RECT 0.587 1.509 0.629 1.551 ;
      RECT 1.119 0.732 1.161 0.774 ;
      RECT 1.195 0.296 1.237 0.338 ;
      RECT 1.195 0.204 1.237 0.246 ;
      RECT 1.195 0.388 1.237 0.43 ;
    LAYER NWELL ;
      RECT -0.115 0.679 2.091 1.773 ;
  END
END AOI22X2_RVT

MACRO AO22X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.744 0.401 0.786 ;
      LAYER M1 ;
        RECT 0.249 0.705 0.404 0.815 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.9 0.553 0.942 ;
      LAYER M1 ;
        RECT 0.401 1.009 0.557 1.119 ;
        RECT 0.507 0.88 0.557 1.009 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.125 0.857 0.167 ;
      LAYER M1 ;
        RECT 0.705 0.097 0.863 0.207 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.6 0.705 0.642 ;
      LAYER M1 ;
        RECT 0.553 0.553 0.708 0.663 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END A4
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.043 0.18 1.085 0.222 ;
        RECT 1.347 0.18 1.389 0.222 ;
        RECT 1.043 0.272 1.085 0.314 ;
        RECT 1.347 0.272 1.389 0.314 ;
        RECT 1.043 0.364 1.085 0.406 ;
        RECT 1.347 0.364 1.389 0.406 ;
        RECT 1.043 0.456 1.085 0.498 ;
        RECT 1.347 0.456 1.389 0.498 ;
        RECT 1.043 0.764 1.085 0.806 ;
        RECT 1.347 0.764 1.389 0.806 ;
        RECT 1.043 0.856 1.085 0.898 ;
        RECT 1.347 0.856 1.389 0.898 ;
        RECT 1.043 0.948 1.085 0.99 ;
        RECT 1.347 0.948 1.389 0.99 ;
        RECT 1.043 1.04 1.085 1.082 ;
        RECT 1.347 1.04 1.389 1.082 ;
        RECT 1.347 1.132 1.389 1.174 ;
        RECT 1.347 1.224 1.389 1.266 ;
        RECT 1.347 1.316 1.389 1.358 ;
        RECT 1.347 1.408 1.389 1.45 ;
      LAYER M1 ;
        RECT 1.344 0.815 1.394 1.47 ;
        RECT 1.039 0.794 1.089 1.102 ;
        RECT 1.313 0.755 1.423 0.815 ;
        RECT 1.011 0.744 1.089 0.794 ;
        RECT 1.313 0.705 1.432 0.755 ;
        RECT 1.011 0.518 1.061 0.744 ;
        RECT 1.382 0.518 1.432 0.705 ;
        RECT 1.011 0.468 1.089 0.518 ;
        RECT 1.344 0.468 1.432 0.518 ;
        RECT 1.039 0.394 1.089 0.468 ;
        RECT 1.344 0.394 1.394 0.468 ;
        RECT 1.039 0.344 1.394 0.394 ;
        RECT 1.039 0.16 1.089 0.344 ;
        RECT 1.344 0.16 1.394 0.344 ;
    END
    ANTENNADIFFAREA 0.2484 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.195 1.298 1.237 1.34 ;
        RECT 1.195 1.39 1.237 1.432 ;
        RECT 0.435 1.407 0.477 1.449 ;
        RECT 1.195 1.482 1.237 1.524 ;
        RECT 0.435 1.499 0.477 1.541 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.672 1.702 ;
        RECT 0.431 1.387 0.481 1.642 ;
        RECT 1.191 1.27 1.241 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.195 0.134 1.237 0.176 ;
        RECT 1.195 0.226 1.237 0.268 ;
        RECT 0.587 0.341 0.629 0.383 ;
      LAYER M1 ;
        RECT 0.583 0.03 0.633 0.403 ;
        RECT 1.191 0.03 1.241 0.288 ;
        RECT 0 -0.03 1.672 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.115 0.568 1.317 0.65 ;
      RECT 0.735 1.152 1.239 1.202 ;
      RECT 1.189 0.65 1.239 1.152 ;
      RECT 0.279 0.503 0.329 0.536 ;
      RECT 0.279 0.27 0.329 0.453 ;
      RECT 0.735 1.202 0.785 1.203 ;
      RECT 0.735 1.029 0.785 1.152 ;
      RECT 0.887 0.503 0.937 1.152 ;
      RECT 0.279 0.453 0.937 0.503 ;
      RECT 0.887 0.27 0.937 0.453 ;
      RECT 0.887 1.337 0.937 1.571 ;
      RECT 0.583 1.337 0.633 1.571 ;
      RECT 0.279 1.287 0.937 1.337 ;
      RECT 0.279 1.337 0.329 1.571 ;
    LAYER PO ;
      RECT 1.429 0.056 1.459 1.597 ;
      RECT 1.277 0.052 1.307 1.604 ;
      RECT 1.581 0.057 1.611 1.598 ;
      RECT 1.125 0.064 1.155 1.604 ;
      RECT 0.213 0.072 0.243 1.621 ;
      RECT 0.821 0.072 0.851 1.621 ;
      RECT 0.973 0.076 1.003 1.621 ;
      RECT 0.061 0.072 0.091 1.621 ;
      RECT 0.365 0.067 0.395 1.621 ;
      RECT 0.517 0.072 0.547 1.621 ;
      RECT 0.669 0.072 0.699 1.621 ;
    LAYER CO ;
      RECT 0.739 1.141 0.781 1.183 ;
      RECT 1.119 0.588 1.161 0.63 ;
      RECT 1.271 0.588 1.313 0.63 ;
      RECT 0.587 1.509 0.629 1.551 ;
      RECT 0.891 0.29 0.933 0.332 ;
      RECT 0.283 1.509 0.325 1.551 ;
      RECT 0.283 1.325 0.325 1.367 ;
      RECT 0.891 1.509 0.933 1.551 ;
      RECT 0.891 1.325 0.933 1.367 ;
      RECT 0.283 0.29 0.325 0.332 ;
      RECT 0.283 0.474 0.325 0.516 ;
      RECT 0.891 0.382 0.933 0.424 ;
      RECT 0.283 1.417 0.325 1.459 ;
      RECT 0.891 0.474 0.933 0.516 ;
      RECT 0.283 0.382 0.325 0.424 ;
      RECT 0.891 1.417 0.933 1.459 ;
      RECT 0.587 1.325 0.629 1.367 ;
      RECT 0.587 1.417 0.629 1.459 ;
      RECT 0.739 1.049 0.781 1.091 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.787 1.773 ;
  END
END AO22X2_RVT

MACRO NOR2X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.665 0.401 0.707 ;
      LAYER M1 ;
        RECT 0.249 0.631 0.421 0.815 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.665 0.553 0.707 ;
      LAYER M1 ;
        RECT 0.489 0.553 0.663 0.733 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.03 ;
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.195 0.151 1.237 0.193 ;
        RECT 1.195 0.245 1.237 0.287 ;
        RECT 1.195 0.337 1.237 0.379 ;
        RECT 1.195 0.43 1.237 0.472 ;
        RECT 1.195 0.841 1.237 0.883 ;
        RECT 1.195 0.933 1.237 0.975 ;
        RECT 1.195 1.027 1.237 1.069 ;
        RECT 1.195 1.119 1.237 1.161 ;
        RECT 1.195 1.212 1.237 1.254 ;
        RECT 1.195 1.304 1.237 1.346 ;
        RECT 1.195 1.398 1.237 1.44 ;
        RECT 1.195 1.49 1.237 1.532 ;
      LAYER M1 ;
        RECT 1.191 0.853 1.241 1.552 ;
        RECT 1.191 0.803 1.551 0.853 ;
        RECT 1.501 0.544 1.551 0.803 ;
        RECT 1.191 0.544 1.241 0.546 ;
        RECT 1.191 0.511 1.551 0.544 ;
        RECT 1.191 0.494 1.575 0.511 ;
        RECT 1.191 0.131 1.241 0.494 ;
        RECT 1.465 0.401 1.575 0.494 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 0.931 0.325 0.973 ;
        RECT 1.347 0.931 1.389 0.973 ;
        RECT 0.739 0.993 0.781 1.035 ;
        RECT 0.283 1.024 0.325 1.066 ;
        RECT 1.043 1.024 1.085 1.066 ;
        RECT 1.347 1.024 1.389 1.066 ;
        RECT 0.739 1.085 0.781 1.127 ;
        RECT 0.283 1.116 0.325 1.158 ;
        RECT 1.043 1.116 1.085 1.158 ;
        RECT 1.347 1.116 1.389 1.158 ;
        RECT 0.283 1.209 0.325 1.251 ;
        RECT 1.043 1.209 1.085 1.251 ;
        RECT 1.347 1.209 1.389 1.251 ;
        RECT 0.283 1.301 0.325 1.343 ;
        RECT 1.043 1.301 1.085 1.343 ;
        RECT 1.347 1.301 1.389 1.343 ;
        RECT 0.283 1.395 0.325 1.437 ;
        RECT 1.043 1.395 1.085 1.437 ;
        RECT 1.347 1.395 1.389 1.437 ;
        RECT 0.283 1.487 0.325 1.529 ;
        RECT 1.043 1.487 1.085 1.529 ;
        RECT 1.347 1.487 1.389 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.672 1.702 ;
        RECT 0.279 0.911 0.329 1.642 ;
        RECT 0.735 0.973 0.785 1.642 ;
        RECT 1.039 1.004 1.089 1.642 ;
        RECT 1.343 0.911 1.393 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.043 0.141 1.085 0.183 ;
        RECT 1.347 0.141 1.389 0.183 ;
        RECT 0.435 0.165 0.477 0.207 ;
        RECT 0.739 0.165 0.781 0.207 ;
        RECT 1.043 0.233 1.085 0.275 ;
        RECT 1.347 0.233 1.389 0.275 ;
        RECT 0.435 0.257 0.477 0.299 ;
        RECT 0.739 0.257 0.781 0.299 ;
        RECT 1.043 0.325 1.085 0.367 ;
        RECT 1.347 0.325 1.389 0.367 ;
      LAYER M1 ;
        RECT 1.039 0.03 1.089 0.387 ;
        RECT 1.343 0.03 1.393 0.387 ;
        RECT 0.431 0.03 0.481 0.319 ;
        RECT 0.735 0.03 0.785 0.319 ;
        RECT 0 -0.03 1.672 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.279 0.383 0.775 0.433 ;
      RECT 0.583 0.802 0.775 0.852 ;
      RECT 0.725 0.666 0.877 0.716 ;
      RECT 0.725 0.433 0.775 0.666 ;
      RECT 0.725 0.716 0.775 0.802 ;
      RECT 0.279 0.131 0.329 0.383 ;
      RECT 0.583 0.131 0.633 0.383 ;
      RECT 0.583 0.852 0.633 1.552 ;
      RECT 1.01 0.661 1.333 0.711 ;
      RECT 0.887 0.501 1.06 0.551 ;
      RECT 0.887 0.803 1.061 0.853 ;
      RECT 1.01 0.551 1.06 0.661 ;
      RECT 1.01 0.711 1.06 0.803 ;
      RECT 0.887 0.853 0.937 1.152 ;
      RECT 0.887 0.792 0.937 0.803 ;
      RECT 0.887 0.131 0.937 0.501 ;
    LAYER PO ;
      RECT 1.125 0.071 1.155 1.612 ;
      RECT 1.277 0.071 1.307 1.612 ;
      RECT 1.429 0.071 1.459 1.612 ;
      RECT 0.821 0.071 0.851 1.612 ;
      RECT 0.973 0.071 1.003 1.612 ;
      RECT 0.061 0.071 0.091 1.612 ;
      RECT 1.581 0.071 1.611 1.612 ;
      RECT 0.213 0.071 0.243 1.612 ;
      RECT 0.669 0.071 0.699 1.612 ;
      RECT 0.365 0.071 0.395 1.612 ;
      RECT 0.517 0.071 0.547 1.612 ;
    LAYER CO ;
      RECT 1.271 0.665 1.313 0.707 ;
      RECT 0.587 0.151 0.629 0.193 ;
      RECT 0.587 0.245 0.629 0.287 ;
      RECT 1.119 0.665 1.161 0.707 ;
      RECT 0.587 1.49 0.629 1.532 ;
      RECT 0.587 1.396 0.629 1.438 ;
      RECT 0.587 1.304 0.629 1.346 ;
      RECT 0.587 1.211 0.629 1.253 ;
      RECT 0.587 0.934 0.629 0.976 ;
      RECT 0.283 0.245 0.325 0.287 ;
      RECT 0.283 0.151 0.325 0.193 ;
      RECT 0.587 1.026 0.629 1.068 ;
      RECT 0.587 1.119 0.629 1.161 ;
      RECT 0.587 0.842 0.629 0.884 ;
      RECT 0.815 0.67 0.857 0.712 ;
      RECT 0.891 0.245 0.933 0.287 ;
      RECT 0.891 0.151 0.933 0.193 ;
      RECT 0.891 0.998 0.933 1.04 ;
      RECT 0.891 0.906 0.933 0.948 ;
      RECT 0.891 0.812 0.933 0.854 ;
      RECT 0.891 1.09 0.933 1.132 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.787 1.773 ;
  END
END NOR2X2_RVT

MACRO NOR4X0_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.665 0.401 0.707 ;
      LAYER M1 ;
        RECT 0.355 0.687 0.405 0.747 ;
        RECT 0.249 0.553 0.405 0.687 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.665 0.553 0.707 ;
      LAYER M1 ;
        RECT 0.401 0.95 0.511 0.967 ;
        RECT 0.401 0.857 0.557 0.95 ;
        RECT 0.507 0.645 0.557 0.857 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.665 0.705 0.707 ;
      LAYER M1 ;
        RECT 0.553 1.007 0.719 1.119 ;
        RECT 0.659 0.645 0.709 1.007 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.665 0.857 0.707 ;
      LAYER M1 ;
        RECT 0.809 0.645 0.967 0.815 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A4
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.499 0.148 1.541 0.19 ;
        RECT 1.499 0.242 1.541 0.284 ;
        RECT 1.499 0.334 1.541 0.376 ;
        RECT 1.499 0.427 1.541 0.469 ;
        RECT 1.499 0.912 1.541 0.954 ;
        RECT 1.499 1.006 1.541 1.048 ;
        RECT 1.499 1.098 1.541 1.14 ;
        RECT 1.499 1.191 1.541 1.233 ;
        RECT 1.499 1.283 1.541 1.325 ;
        RECT 1.499 1.377 1.541 1.419 ;
        RECT 1.499 1.469 1.541 1.511 ;
      LAYER M1 ;
        RECT 1.495 0.942 1.545 1.531 ;
        RECT 1.495 0.892 1.699 0.942 ;
        RECT 1.649 0.511 1.699 0.892 ;
        RECT 1.617 0.487 1.727 0.511 ;
        RECT 1.495 0.487 1.545 0.489 ;
        RECT 1.495 0.437 1.727 0.487 ;
        RECT 1.495 0.128 1.545 0.437 ;
        RECT 1.617 0.401 1.727 0.437 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 0.93 0.325 0.972 ;
        RECT 1.347 1.021 1.389 1.063 ;
        RECT 0.283 1.024 0.325 1.066 ;
        RECT 1.043 1.074 1.085 1.116 ;
        RECT 1.347 1.113 1.389 1.155 ;
        RECT 0.283 1.116 0.325 1.158 ;
        RECT 1.043 1.166 1.085 1.208 ;
        RECT 1.347 1.206 1.389 1.248 ;
        RECT 0.283 1.209 0.325 1.251 ;
        RECT 1.347 1.298 1.389 1.34 ;
        RECT 0.283 1.301 0.325 1.343 ;
        RECT 1.347 1.392 1.389 1.434 ;
        RECT 0.283 1.395 0.325 1.437 ;
        RECT 1.347 1.484 1.389 1.526 ;
        RECT 0.283 1.487 0.325 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.824 1.702 ;
        RECT 0.279 0.91 0.329 1.642 ;
        RECT 1.039 1.054 1.089 1.642 ;
        RECT 1.343 1.001 1.393 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.043 0.138 1.085 0.18 ;
        RECT 1.347 0.138 1.389 0.18 ;
        RECT 1.043 0.23 1.085 0.272 ;
        RECT 1.347 0.23 1.389 0.272 ;
        RECT 0.435 0.269 0.477 0.311 ;
        RECT 0.739 0.28 0.781 0.322 ;
        RECT 1.347 0.322 1.389 0.364 ;
      LAYER M1 ;
        RECT 1.343 0.03 1.393 0.384 ;
        RECT 0.735 0.03 0.785 0.342 ;
        RECT 0.431 0.03 0.481 0.331 ;
        RECT 1.039 0.03 1.089 0.292 ;
        RECT 0 -0.03 1.824 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.279 0.397 1.083 0.447 ;
      RECT 0.887 0.903 1.083 0.953 ;
      RECT 1.033 0.747 1.181 0.797 ;
      RECT 1.033 0.447 1.083 0.747 ;
      RECT 1.033 0.797 1.083 0.903 ;
      RECT 0.279 0.261 0.329 0.397 ;
      RECT 0.583 0.261 0.633 0.397 ;
      RECT 0.887 0.26 0.937 0.397 ;
      RECT 0.887 0.953 0.937 1.535 ;
      RECT 0.887 0.883 0.937 0.903 ;
      RECT 1.191 0.498 1.365 0.548 ;
      RECT 1.192 0.85 1.365 0.875 ;
      RECT 1.191 0.875 1.365 0.9 ;
      RECT 1.314 0.661 1.485 0.711 ;
      RECT 1.314 0.548 1.364 0.661 ;
      RECT 1.314 0.711 1.364 0.85 ;
      RECT 1.191 0.128 1.241 0.498 ;
      RECT 1.191 0.9 1.241 1.224 ;
    LAYER PO ;
      RECT 1.429 0.068 1.459 1.609 ;
      RECT 1.581 0.068 1.611 1.609 ;
      RECT 1.125 0.068 1.155 1.609 ;
      RECT 1.277 0.068 1.307 1.609 ;
      RECT 0.973 0.068 1.003 1.609 ;
      RECT 1.733 0.072 1.763 1.609 ;
      RECT 0.061 0.072 0.091 1.609 ;
      RECT 0.821 0.072 0.851 1.609 ;
      RECT 0.213 0.072 0.243 1.609 ;
      RECT 0.669 0.072 0.699 1.609 ;
      RECT 0.365 0.072 0.395 1.609 ;
      RECT 0.517 0.072 0.547 1.609 ;
    LAYER CO ;
      RECT 0.891 1.458 0.933 1.5 ;
      RECT 0.891 1.366 0.933 1.408 ;
      RECT 0.891 1.272 0.933 1.314 ;
      RECT 0.891 1.18 0.933 1.222 ;
      RECT 1.423 0.665 1.465 0.707 ;
      RECT 1.195 1.162 1.237 1.204 ;
      RECT 1.195 0.978 1.237 1.02 ;
      RECT 0.891 1.087 0.933 1.129 ;
      RECT 0.587 0.281 0.629 0.323 ;
      RECT 0.891 0.903 0.933 0.945 ;
      RECT 1.195 0.884 1.237 0.926 ;
      RECT 1.195 1.07 1.237 1.112 ;
      RECT 0.891 0.995 0.933 1.037 ;
      RECT 1.119 0.751 1.161 0.793 ;
      RECT 1.195 0.242 1.237 0.284 ;
      RECT 1.195 0.148 1.237 0.19 ;
      RECT 0.891 0.28 0.933 0.322 ;
      RECT 0.283 0.281 0.325 0.323 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.939 1.773 ;
  END
END NOR4X0_RVT

MACRO AND4X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.28 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 1.043 0.857 1.085 ;
      LAYER M1 ;
        RECT 0.705 1.089 0.815 1.119 ;
        RECT 0.705 1.039 0.877 1.089 ;
        RECT 0.705 1.009 0.815 1.039 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0165 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.739 0.705 0.781 ;
      LAYER M1 ;
        RECT 0.553 0.785 0.663 0.815 ;
        RECT 0.553 0.735 0.725 0.785 ;
        RECT 0.553 0.705 0.663 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0165 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.043 0.553 1.085 ;
      LAYER M1 ;
        RECT 0.401 1.089 0.511 1.119 ;
        RECT 0.401 1.039 0.573 1.089 ;
        RECT 0.401 1.009 0.511 1.039 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0165 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.249 0.785 0.359 0.815 ;
        RECT 0.249 0.735 0.421 0.785 ;
        RECT 0.249 0.705 0.359 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0165 ;
  END A4
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.803 0.148 1.845 0.19 ;
        RECT 1.803 0.24 1.845 0.282 ;
        RECT 1.803 0.332 1.845 0.374 ;
        RECT 1.803 0.424 1.845 0.466 ;
        RECT 1.803 0.935 1.845 0.977 ;
        RECT 1.803 1.027 1.845 1.069 ;
        RECT 1.803 1.119 1.845 1.161 ;
        RECT 1.803 1.211 1.845 1.253 ;
        RECT 1.803 1.303 1.845 1.345 ;
        RECT 1.803 1.395 1.845 1.437 ;
        RECT 1.803 1.487 1.845 1.529 ;
      LAYER M1 ;
        RECT 1.799 0.793 1.849 1.564 ;
        RECT 1.799 0.743 2.094 0.793 ;
        RECT 2.044 0.663 2.094 0.743 ;
        RECT 2.044 0.59 2.183 0.663 ;
        RECT 1.799 0.553 2.183 0.59 ;
        RECT 1.799 0.54 2.094 0.553 ;
        RECT 1.799 0.12 1.849 0.54 ;
    END
    ANTENNADIFFAREA 0.1488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.651 0.843 1.693 0.885 ;
        RECT 1.651 0.935 1.693 0.977 ;
        RECT 1.955 0.935 1.997 0.977 ;
        RECT 1.651 1.027 1.693 1.069 ;
        RECT 1.955 1.027 1.997 1.069 ;
        RECT 1.347 1.119 1.389 1.161 ;
        RECT 1.651 1.119 1.693 1.161 ;
        RECT 1.955 1.119 1.997 1.161 ;
        RECT 1.347 1.211 1.389 1.253 ;
        RECT 1.651 1.211 1.693 1.253 ;
        RECT 1.955 1.211 1.997 1.253 ;
        RECT 1.043 1.219 1.085 1.261 ;
        RECT 1.347 1.303 1.389 1.345 ;
        RECT 1.651 1.303 1.693 1.345 ;
        RECT 1.955 1.303 1.997 1.345 ;
        RECT 1.043 1.311 1.085 1.353 ;
        RECT 1.347 1.395 1.389 1.437 ;
        RECT 1.651 1.395 1.693 1.437 ;
        RECT 1.955 1.395 1.997 1.437 ;
        RECT 1.043 1.403 1.085 1.445 ;
        RECT 0.435 1.405 0.477 1.447 ;
        RECT 0.739 1.405 0.781 1.447 ;
        RECT 1.347 1.487 1.389 1.529 ;
        RECT 1.651 1.487 1.693 1.529 ;
        RECT 1.955 1.487 1.997 1.529 ;
        RECT 1.043 1.495 1.085 1.537 ;
        RECT 0.435 1.497 0.477 1.539 ;
        RECT 0.739 1.497 0.781 1.539 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 2.28 1.702 ;
        RECT 0.431 1.385 0.481 1.642 ;
        RECT 0.735 1.385 0.785 1.642 ;
        RECT 1.039 1.199 1.089 1.642 ;
        RECT 1.343 1.099 1.393 1.642 ;
        RECT 1.647 0.823 1.697 1.642 ;
        RECT 1.951 0.915 2.001 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 0.283 0.141 0.325 0.183 ;
        RECT 1.347 0.148 1.389 0.19 ;
        RECT 1.651 0.148 1.693 0.19 ;
        RECT 1.955 0.148 1.997 0.19 ;
        RECT 1.043 0.15 1.085 0.192 ;
        RECT 0.283 0.233 0.325 0.275 ;
        RECT 1.347 0.24 1.389 0.282 ;
        RECT 1.651 0.24 1.693 0.282 ;
        RECT 1.955 0.24 1.997 0.282 ;
        RECT 1.043 0.242 1.085 0.284 ;
        RECT 0.283 0.325 0.325 0.367 ;
        RECT 1.651 0.332 1.693 0.374 ;
        RECT 1.955 0.332 1.997 0.374 ;
        RECT 0.283 0.417 0.325 0.459 ;
        RECT 1.651 0.424 1.693 0.466 ;
        RECT 1.955 0.424 1.997 0.466 ;
      LAYER M1 ;
        RECT 1.647 0.03 1.697 0.486 ;
        RECT 1.951 0.03 2.001 0.486 ;
        RECT 0.279 0.03 0.329 0.479 ;
        RECT 1.039 0.03 1.089 0.304 ;
        RECT 1.343 0.03 1.393 0.302 ;
        RECT 0 -0.03 2.28 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.891 0.325 0.933 0.367 ;
      RECT 0.891 0.417 0.933 0.459 ;
      RECT 1.195 0.15 1.237 0.192 ;
      RECT 1.119 0.66 1.161 0.702 ;
      RECT 1.195 0.242 1.237 0.284 ;
      RECT 0.891 1.497 0.933 1.539 ;
      RECT 1.499 1.211 1.541 1.253 ;
      RECT 1.195 1.219 1.237 1.261 ;
      RECT 0.283 1.405 0.325 1.447 ;
      RECT 1.195 0.15 1.237 0.192 ;
      RECT 0.283 1.497 0.325 1.539 ;
      RECT 1.499 1.303 1.541 1.345 ;
      RECT 0.891 0.141 0.933 0.183 ;
      RECT 1.423 0.733 1.465 0.775 ;
      RECT 1.499 0.148 1.541 0.19 ;
      RECT 1.879 0.644 1.921 0.686 ;
      RECT 1.727 0.644 1.769 0.686 ;
      RECT 1.195 1.311 1.237 1.353 ;
      RECT 1.195 1.495 1.237 1.537 ;
      RECT 1.195 1.311 1.237 1.353 ;
      RECT 0.587 1.405 0.629 1.447 ;
      RECT 0.587 1.497 0.629 1.539 ;
      RECT 1.499 1.487 1.541 1.529 ;
      RECT 1.195 1.495 1.237 1.537 ;
      RECT 1.499 0.24 1.541 0.282 ;
      RECT 1.499 0.148 1.541 0.19 ;
      RECT 1.499 1.395 1.541 1.437 ;
      RECT 1.499 1.395 1.541 1.437 ;
      RECT 1.499 1.303 1.541 1.345 ;
      RECT 0.891 1.405 0.933 1.447 ;
      RECT 1.499 1.119 1.541 1.161 ;
      RECT 1.195 1.403 1.237 1.445 ;
      RECT 1.195 1.403 1.237 1.445 ;
      RECT 1.195 1.219 1.237 1.261 ;
      RECT 0.891 0.233 0.933 0.275 ;
      RECT 1.499 1.487 1.541 1.529 ;
      RECT 1.499 1.211 1.541 1.253 ;
    LAYER M1 ;
      RECT 1.535 0.64 1.941 0.69 ;
      RECT 1.495 1.071 1.545 1.564 ;
      RECT 1.495 1.021 1.585 1.071 ;
      RECT 1.495 0.12 1.545 0.461 ;
      RECT 1.495 0.461 1.585 0.511 ;
      RECT 1.535 0.511 1.585 0.64 ;
      RECT 1.535 0.69 1.585 1.021 ;
      RECT 0.927 0.672 1.181 0.706 ;
      RECT 0.887 0.656 1.181 0.672 ;
      RECT 0.279 1.313 0.329 1.559 ;
      RECT 0.583 1.313 0.633 1.559 ;
      RECT 0.279 1.263 0.977 1.313 ;
      RECT 0.887 0.121 0.937 0.622 ;
      RECT 0.887 1.313 0.937 1.559 ;
      RECT 0.927 0.706 0.977 1.263 ;
      RECT 0.887 0.622 0.977 0.656 ;
      RECT 1.29 0.729 1.485 0.779 ;
      RECT 1.191 0.99 1.241 1.557 ;
      RECT 1.191 0.94 1.34 0.99 ;
      RECT 1.191 0.117 1.241 0.551 ;
      RECT 1.191 0.551 1.315 0.553 ;
      RECT 1.191 0.553 1.34 0.601 ;
      RECT 1.29 0.779 1.34 0.94 ;
      RECT 1.29 0.601 1.34 0.729 ;
    LAYER PO ;
      RECT 1.277 0.072 1.307 1.609 ;
      RECT 1.429 0.062 1.459 1.609 ;
      RECT 1.125 0.072 1.155 1.609 ;
      RECT 0.973 0.071 1.003 1.609 ;
      RECT 0.669 0.071 0.699 1.609 ;
      RECT 0.365 0.071 0.395 1.609 ;
      RECT 0.517 0.071 0.547 1.609 ;
      RECT 0.213 0.071 0.243 1.609 ;
      RECT 0.821 0.071 0.851 1.609 ;
      RECT 0.061 0.071 0.091 1.609 ;
      RECT 1.733 0.062 1.763 1.609 ;
      RECT 1.885 0.062 1.915 1.609 ;
      RECT 2.189 0.062 2.219 1.609 ;
      RECT 2.037 0.062 2.067 1.609 ;
      RECT 1.581 0.062 1.611 1.609 ;
    LAYER NWELL ;
      RECT -0.115 0.679 2.395 1.773 ;
  END
END AND4X2_RVT

MACRO MUX41X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 3.344 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.727 0.133 1.769 0.175 ;
      LAYER M1 ;
        RECT 1.707 0.097 1.879 0.207 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A1
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.967 0.814 1.009 0.856 ;
      LAYER M1 ;
        RECT 0.857 0.86 0.967 0.967 ;
        RECT 0.857 0.81 1.037 0.86 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A3
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.575 0.748 1.617 0.79 ;
      LAYER M1 ;
        RECT 1.465 0.699 1.637 0.822 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A2
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.623 0.857 0.665 ;
      LAYER M1 ;
        RECT 0.812 0.553 0.967 0.685 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A4
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 2.183 1.448 2.225 1.49 ;
        RECT 2.639 1.448 2.681 1.49 ;
      LAYER M1 ;
        RECT 2.529 1.494 2.659 1.581 ;
        RECT 2.162 1.444 2.708 1.494 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.09 0.553 0.132 ;
        RECT 0.663 0.09 0.705 0.132 ;
        RECT 1.271 0.09 1.313 0.132 ;
        RECT 1.423 0.092 1.465 0.134 ;
        RECT 0.359 0.126 0.401 0.168 ;
      LAYER M1 ;
        RECT 0.659 0.278 1.14 0.328 ;
        RECT 0.659 0.138 0.709 0.278 ;
        RECT 1.09 0.138 1.14 0.278 ;
        RECT 0.249 0.138 0.417 0.207 ;
        RECT 0.249 0.088 0.725 0.138 ;
        RECT 1.09 0.088 1.485 0.138 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.072 ;
  END S1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 3.019 0.276 3.061 0.318 ;
        RECT 3.019 0.368 3.061 0.41 ;
        RECT 3.019 0.969 3.061 1.011 ;
        RECT 3.019 1.061 3.061 1.103 ;
      LAYER M1 ;
        RECT 3.015 0.971 3.065 1.146 ;
        RECT 3.015 0.921 3.19 0.971 ;
        RECT 3.14 0.768 3.19 0.921 ;
        RECT 3.137 0.553 3.248 0.768 ;
        RECT 3.14 0.453 3.19 0.553 ;
        RECT 3.015 0.403 3.19 0.453 ;
        RECT 3.015 0.216 3.065 0.403 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.073 0.325 1.115 ;
        RECT 0.283 1.165 0.325 1.207 ;
        RECT 2.563 1.212 2.605 1.254 ;
        RECT 1.651 1.32 1.693 1.362 ;
        RECT 0.891 1.344 0.933 1.386 ;
        RECT 2.867 1.412 2.909 1.454 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
        RECT 2.639 1.651 2.681 1.693 ;
        RECT 2.791 1.651 2.833 1.693 ;
        RECT 2.943 1.651 2.985 1.693 ;
        RECT 3.095 1.651 3.137 1.693 ;
        RECT 3.247 1.651 3.289 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 3.344 1.702 ;
        RECT 3.097 1.488 3.147 1.642 ;
        RECT 0.887 1.324 0.937 1.642 ;
        RECT 1.647 1.3 1.697 1.642 ;
        RECT 2.863 1.438 3.147 1.488 ;
        RECT 0.279 1.05 0.329 1.642 ;
        RECT 2.863 1.258 2.913 1.438 ;
        RECT 2.543 1.208 2.913 1.258 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 2.639 -0.021 2.681 0.021 ;
        RECT 2.791 -0.021 2.833 0.021 ;
        RECT 2.943 -0.021 2.985 0.021 ;
        RECT 3.095 -0.021 3.137 0.021 ;
        RECT 3.247 -0.021 3.289 0.021 ;
        RECT 2.867 0.159 2.909 0.201 ;
        RECT 0.891 0.182 0.933 0.224 ;
        RECT 2.563 0.196 2.605 0.238 ;
        RECT 1.651 0.261 1.693 0.303 ;
        RECT 0.283 0.461 0.325 0.503 ;
        RECT 0.283 0.553 0.325 0.595 ;
      LAYER M1 ;
        RECT 0.279 0.462 0.329 0.625 ;
        RECT 0.131 0.412 0.329 0.462 ;
        RECT 1.535 0.257 1.713 0.307 ;
        RECT 2.543 0.192 2.801 0.242 ;
        RECT 0.867 0.178 0.978 0.228 ;
        RECT 0.131 0.03 0.181 0.412 ;
        RECT 1.535 0.03 1.585 0.257 ;
        RECT 2.863 0.03 2.913 0.223 ;
        RECT 2.751 0.03 2.801 0.192 ;
        RECT 0.928 0.03 0.978 0.178 ;
        RECT 0 -0.03 3.344 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.511 1.537 0.553 1.579 ;
      RECT 2.107 0.818 2.149 0.86 ;
      RECT 1.271 1.538 1.313 1.58 ;
      RECT 2.183 0.092 2.225 0.134 ;
      RECT 1.955 0.915 1.997 0.957 ;
      RECT 1.119 0.587 1.161 0.629 ;
      RECT 0.435 1.073 0.477 1.115 ;
      RECT 1.879 0.8 1.921 0.842 ;
      RECT 2.335 1.348 2.377 1.39 ;
      RECT 2.639 0.09 2.681 0.132 ;
      RECT 0.587 0.404 0.629 0.446 ;
      RECT 2.411 0.818 2.453 0.86 ;
      RECT 0.587 1.322 0.629 1.364 ;
      RECT 1.195 1.038 1.237 1.08 ;
      RECT 2.715 0.798 2.757 0.84 ;
      RECT 2.715 0.412 2.757 0.454 ;
      RECT 0.435 1.165 0.477 1.207 ;
      RECT 2.031 0.092 2.073 0.134 ;
      RECT 2.259 0.512 2.301 0.554 ;
      RECT 2.259 0.818 2.301 0.86 ;
      RECT 0.435 1.257 0.477 1.299 ;
      RECT 0.435 0.492 0.477 0.534 ;
      RECT 2.943 0.662 2.985 0.704 ;
      RECT 2.031 1.432 2.073 1.474 ;
      RECT 2.411 0.512 2.453 0.554 ;
      RECT 2.335 0.092 2.377 0.134 ;
      RECT 1.347 0.481 1.389 0.523 ;
      RECT 0.663 1.439 0.705 1.481 ;
      RECT 1.347 1.248 1.389 1.29 ;
      RECT 1.879 0.657 1.921 0.699 ;
      RECT 1.423 1.422 1.465 1.464 ;
      RECT 1.119 1.504 1.161 1.546 ;
      RECT 1.955 0.462 1.997 0.504 ;
      RECT 1.195 0.383 1.237 0.425 ;
      RECT 2.107 0.512 2.149 0.554 ;
    LAYER M1 ;
      RECT 1.443 1.1 1.753 1.15 ;
      RECT 1.703 0.736 1.753 1.1 ;
      RECT 1.856 0.652 1.941 0.686 ;
      RECT 1.703 0.702 1.906 0.736 ;
      RECT 1.703 0.686 1.941 0.702 ;
      RECT 0.431 1.434 0.733 1.484 ;
      RECT 0.683 1.174 0.733 1.434 ;
      RECT 0.431 0.472 0.481 1.434 ;
      RECT 1.419 1.426 1.469 1.484 ;
      RECT 1.115 1.376 1.493 1.426 ;
      RECT 1.443 1.15 1.493 1.376 ;
      RECT 1.069 0.934 1.165 0.984 ;
      RECT 1.115 1.184 1.165 1.376 ;
      RECT 1.069 1.174 1.165 1.184 ;
      RECT 1.069 0.984 1.119 1.124 ;
      RECT 0.683 1.134 1.165 1.174 ;
      RECT 1.115 0.557 1.165 0.934 ;
      RECT 0.683 1.124 1.119 1.134 ;
      RECT 1.935 0.911 2.045 0.961 ;
      RECT 1.343 0.458 2.153 0.508 ;
      RECT 1.995 0.508 2.045 0.911 ;
      RECT 2.103 0.508 2.153 0.88 ;
      RECT 1.343 0.508 1.393 1.31 ;
      RECT 2.401 1.104 2.761 1.154 ;
      RECT 2.711 0.392 2.761 1.104 ;
      RECT 2.401 1.154 2.451 1.344 ;
      RECT 2.056 1.344 2.451 1.394 ;
      RECT 2.009 1.428 2.106 1.478 ;
      RECT 2.056 1.394 2.106 1.428 ;
      RECT 2.255 0.933 2.634 0.983 ;
      RECT 2.584 0.342 2.634 0.933 ;
      RECT 2.584 0.292 2.928 0.342 ;
      RECT 2.878 0.342 2.928 0.658 ;
      RECT 2.878 0.658 3.005 0.708 ;
      RECT 2.255 0.492 2.305 0.933 ;
      RECT 1.115 1.526 1.165 1.578 ;
      RECT 0.987 1.476 1.165 1.526 ;
      RECT 0.987 1.274 1.037 1.476 ;
      RECT 0.783 1.224 1.037 1.274 ;
      RECT 0.483 1.534 0.833 1.584 ;
      RECT 0.783 1.274 0.833 1.534 ;
      RECT 2.407 0.407 2.457 0.88 ;
      RECT 1.219 0.357 2.457 0.378 ;
      RECT 0.583 0.378 2.457 0.407 ;
      RECT 0.583 0.428 0.633 1.384 ;
      RECT 1.169 1.034 1.269 1.084 ;
      RECT 0.583 0.407 1.269 0.428 ;
      RECT 1.219 0.428 1.269 1.034 ;
      RECT 1.547 1.2 1.853 1.25 ;
      RECT 1.803 0.796 1.941 0.846 ;
      RECT 1.803 0.846 1.853 1.2 ;
      RECT 1.245 1.534 1.597 1.584 ;
      RECT 1.547 1.25 1.597 1.534 ;
      RECT 2.004 0.088 2.245 0.138 ;
      RECT 2.315 0.088 2.701 0.138 ;
    LAYER PO ;
      RECT 1.581 0.071 1.611 1.609 ;
      RECT 1.733 0.071 1.763 1.609 ;
      RECT 2.189 0.748 2.219 1.609 ;
      RECT 2.189 0.069 2.219 0.648 ;
      RECT 1.429 0.071 1.459 0.673 ;
      RECT 1.429 0.821 1.459 1.609 ;
      RECT 0.517 0.071 0.547 1.609 ;
      RECT 0.213 0.071 0.243 1.609 ;
      RECT 3.101 0.072 3.131 1.61 ;
      RECT 0.973 0.071 1.003 1.609 ;
      RECT 2.645 0.072 2.675 1.61 ;
      RECT 1.885 0.071 1.915 0.7 ;
      RECT 1.885 0.8 1.915 1.609 ;
      RECT 2.341 0.069 2.371 0.624 ;
      RECT 2.797 0.072 2.827 1.61 ;
      RECT 1.125 0.071 1.155 0.627 ;
      RECT 1.277 0.072 1.307 1.61 ;
      RECT 1.125 0.756 1.155 1.609 ;
      RECT 0.669 0.071 0.699 0.627 ;
      RECT 3.253 0.072 3.283 1.61 ;
      RECT 0.061 0.071 0.091 1.609 ;
      RECT 2.037 0.069 2.067 1.609 ;
      RECT 0.669 0.75 0.699 1.609 ;
      RECT 0.365 0.071 0.395 1.609 ;
      RECT 2.949 0.072 2.979 1.61 ;
      RECT 2.341 0.748 2.371 1.609 ;
      RECT 0.821 0.071 0.851 1.609 ;
      RECT 2.493 0.071 2.523 1.609 ;
    LAYER NWELL ;
      RECT -0.115 0.679 3.459 1.773 ;
  END
END MUX41X1_RVT

MACRO OA21X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.672 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.271 0.814 0.421 0.817 ;
        RECT 0.249 0.717 0.421 0.814 ;
        RECT 0.249 0.705 0.359 0.717 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.027 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.482 0.553 1.524 ;
      LAYER M1 ;
        RECT 0.401 1.571 0.511 1.575 ;
        RECT 0.401 1.465 0.573 1.571 ;
        RECT 0.426 1.46 0.573 1.465 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.027 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.827 0.857 0.869 ;
      LAYER M1 ;
        RECT 0.712 0.962 0.861 0.986 ;
        RECT 0.705 0.853 0.861 0.962 ;
        RECT 0.811 0.807 0.861 0.853 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0132 ;
  END A3
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.043 0.239 1.085 0.281 ;
        RECT 1.347 0.239 1.389 0.281 ;
        RECT 1.043 0.331 1.085 0.373 ;
        RECT 1.347 0.331 1.389 0.373 ;
        RECT 1.043 0.423 1.085 0.465 ;
        RECT 1.347 0.423 1.389 0.465 ;
        RECT 1.043 0.987 1.085 1.029 ;
        RECT 1.347 0.987 1.389 1.029 ;
        RECT 1.043 1.079 1.085 1.121 ;
        RECT 1.347 1.079 1.389 1.121 ;
        RECT 1.043 1.171 1.085 1.213 ;
        RECT 1.347 1.171 1.389 1.213 ;
        RECT 1.043 1.263 1.085 1.305 ;
        RECT 1.347 1.263 1.389 1.305 ;
        RECT 1.043 1.355 1.085 1.397 ;
        RECT 1.347 1.355 1.389 1.397 ;
      LAYER M1 ;
        RECT 1.039 1.006 1.089 1.426 ;
        RECT 1.343 1.006 1.393 1.426 ;
        RECT 1.039 0.956 1.532 1.006 ;
        RECT 1.482 0.542 1.532 0.956 ;
        RECT 1.039 0.53 1.532 0.542 ;
        RECT 1.039 0.492 1.591 0.53 ;
        RECT 1.039 0.188 1.089 0.492 ;
        RECT 1.343 0.188 1.393 0.492 ;
        RECT 1.455 0.392 1.591 0.492 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 0.987 0.325 1.029 ;
        RECT 0.283 1.079 0.325 1.121 ;
        RECT 0.283 1.171 0.325 1.213 ;
        RECT 1.195 1.171 1.237 1.213 ;
        RECT 0.283 1.263 0.325 1.305 ;
        RECT 0.891 1.263 0.933 1.305 ;
        RECT 1.195 1.263 1.237 1.305 ;
        RECT 0.283 1.355 0.325 1.397 ;
        RECT 0.891 1.355 0.933 1.397 ;
        RECT 1.195 1.355 1.237 1.397 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.672 1.702 ;
        RECT 0.279 0.958 0.329 1.642 ;
        RECT 0.887 1.243 0.937 1.642 ;
        RECT 1.191 1.133 1.241 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.195 0.203 1.237 0.245 ;
        RECT 0.435 0.239 0.477 0.281 ;
        RECT 1.195 0.295 1.237 0.337 ;
        RECT 0.435 0.331 0.477 0.373 ;
        RECT 0.435 0.423 0.477 0.465 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.512 ;
        RECT 1.191 0.03 1.241 0.399 ;
        RECT 0 -0.03 1.672 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.231 0.681 1.317 0.699 ;
      RECT 1.231 0.613 1.317 0.631 ;
      RECT 0.887 0.631 1.317 0.681 ;
      RECT 0.583 1.18 0.633 1.393 ;
      RECT 0.583 1.106 0.633 1.13 ;
      RECT 0.735 1.18 0.785 1.393 ;
      RECT 0.735 1.106 0.785 1.13 ;
      RECT 1.07 0.681 1.156 0.699 ;
      RECT 1.07 0.613 1.156 0.631 ;
      RECT 0.913 0.681 0.963 1.13 ;
      RECT 0.887 0.181 0.937 0.631 ;
      RECT 0.583 1.13 0.963 1.18 ;
      RECT 0.279 0.598 0.633 0.648 ;
      RECT 0.735 0.181 0.785 0.412 ;
      RECT 0.583 0.412 0.785 0.462 ;
      RECT 0.583 0.462 0.633 0.598 ;
      RECT 0.583 0.181 0.633 0.412 ;
      RECT 0.279 0.178 0.329 0.598 ;
    LAYER PO ;
      RECT 0.973 0.101 1.003 1.469 ;
      RECT 1.125 0.069 1.155 1.608 ;
      RECT 0.365 0.101 0.395 1.469 ;
      RECT 0.821 0.101 0.851 1.469 ;
      RECT 1.429 0.101 1.459 1.469 ;
      RECT 1.581 0.101 1.611 1.469 ;
      RECT 0.061 0.101 0.091 1.469 ;
      RECT 1.277 0.069 1.307 1.608 ;
      RECT 0.517 0.101 0.547 1.567 ;
      RECT 0.213 0.101 0.243 1.469 ;
      RECT 0.669 0.101 0.699 1.469 ;
    LAYER CO ;
      RECT 0.587 0.331 0.629 0.373 ;
      RECT 1.271 0.635 1.313 0.677 ;
      RECT 0.891 0.211 0.933 0.253 ;
      RECT 0.891 0.303 0.933 0.345 ;
      RECT 0.283 0.239 0.325 0.281 ;
      RECT 0.739 1.23 0.781 1.272 ;
      RECT 0.739 1.322 0.781 1.364 ;
      RECT 0.587 0.423 0.629 0.465 ;
      RECT 0.283 0.423 0.325 0.465 ;
      RECT 0.283 0.331 0.325 0.373 ;
      RECT 0.739 0.303 0.781 0.345 ;
      RECT 0.739 0.211 0.781 0.253 ;
      RECT 0.587 1.23 0.629 1.272 ;
      RECT 0.587 1.322 0.629 1.364 ;
      RECT 1.119 0.635 1.161 0.677 ;
      RECT 0.587 1.138 0.629 1.18 ;
      RECT 0.587 0.239 0.629 0.281 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.787 1.787 ;
  END
END OA21X2_RVT

MACRO OA221X2_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.976 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.739 0.401 0.781 ;
      LAYER M1 ;
        RECT 0.271 0.81 0.421 0.817 ;
        RECT 0.249 0.71 0.421 0.81 ;
        RECT 0.249 0.701 0.359 0.71 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.482 0.553 1.524 ;
      LAYER M1 ;
        RECT 0.401 1.571 0.511 1.577 ;
        RECT 0.401 1.461 0.573 1.571 ;
        RECT 0.426 1.46 0.573 1.461 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.866 0.857 0.908 ;
      LAYER M1 ;
        RECT 0.811 1.002 0.968 1.139 ;
        RECT 0.811 0.842 0.861 1.002 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.739 0.705 0.781 ;
      LAYER M1 ;
        RECT 0.56 0.963 0.709 0.986 ;
        RECT 0.553 0.854 0.709 0.963 ;
        RECT 0.659 0.713 0.709 0.854 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.119 0.739 1.161 0.781 ;
      LAYER M1 ;
        RECT 1.115 0.675 1.165 0.808 ;
        RECT 1.023 0.658 1.165 0.675 ;
        RECT 1.009 0.601 1.165 0.658 ;
        RECT 1.009 0.549 1.123 0.601 ;
        RECT 1.023 0.541 1.123 0.549 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0177 ;
  END A5
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.347 0.239 1.389 0.281 ;
        RECT 1.651 0.239 1.693 0.281 ;
        RECT 1.347 0.331 1.389 0.373 ;
        RECT 1.651 0.331 1.693 0.373 ;
        RECT 1.347 0.423 1.389 0.465 ;
        RECT 1.651 0.423 1.693 0.465 ;
        RECT 1.347 0.987 1.389 1.029 ;
        RECT 1.651 0.987 1.693 1.029 ;
        RECT 1.347 1.079 1.389 1.121 ;
        RECT 1.651 1.079 1.693 1.121 ;
        RECT 1.347 1.171 1.389 1.213 ;
        RECT 1.651 1.171 1.693 1.213 ;
        RECT 1.347 1.263 1.389 1.305 ;
        RECT 1.651 1.263 1.693 1.305 ;
        RECT 1.347 1.355 1.389 1.397 ;
        RECT 1.651 1.355 1.693 1.397 ;
      LAYER M1 ;
        RECT 1.343 1.006 1.393 1.426 ;
        RECT 1.647 1.006 1.697 1.426 ;
        RECT 1.343 0.956 1.836 1.006 ;
        RECT 1.786 0.542 1.836 0.956 ;
        RECT 1.343 0.53 1.836 0.542 ;
        RECT 1.343 0.492 1.911 0.53 ;
        RECT 1.343 0.188 1.393 0.492 ;
        RECT 1.647 0.188 1.697 0.492 ;
        RECT 1.751 0.392 1.911 0.492 ;
    END
    ANTENNADIFFAREA 0.2488 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 1.079 0.325 1.121 ;
        RECT 0.283 1.171 0.325 1.213 ;
        RECT 1.499 1.171 1.541 1.213 ;
        RECT 0.283 1.263 0.325 1.305 ;
        RECT 1.499 1.263 1.541 1.305 ;
        RECT 0.283 1.355 0.325 1.397 ;
        RECT 0.891 1.355 0.933 1.397 ;
        RECT 1.043 1.355 1.085 1.397 ;
        RECT 1.499 1.355 1.541 1.397 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.976 1.702 ;
        RECT 0.279 0.958 0.329 1.642 ;
        RECT 0.887 1.335 0.937 1.642 ;
        RECT 1.039 1.333 1.089 1.642 ;
        RECT 1.495 1.133 1.545 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 1.499 0.203 1.541 0.245 ;
        RECT 0.435 0.239 0.477 0.281 ;
        RECT 1.499 0.295 1.541 0.337 ;
        RECT 0.435 0.331 0.477 0.373 ;
        RECT 0.435 0.423 0.477 0.465 ;
      LAYER M1 ;
        RECT 0.431 0.03 0.481 0.512 ;
        RECT 1.495 0.03 1.545 0.399 ;
        RECT 0 -0.03 1.976 0.03 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.535 0.681 1.621 0.699 ;
      RECT 1.535 0.613 1.621 0.631 ;
      RECT 1.227 0.631 1.621 0.681 ;
      RECT 0.583 1.263 0.633 1.393 ;
      RECT 0.583 1.106 0.633 1.213 ;
      RECT 1.383 0.681 1.469 0.699 ;
      RECT 1.383 0.613 1.469 0.631 ;
      RECT 1.191 0.483 1.277 0.533 ;
      RECT 1.039 0.903 1.277 0.953 ;
      RECT 1.227 0.533 1.277 0.631 ;
      RECT 1.191 0.211 1.241 0.483 ;
      RECT 1.191 0.953 1.241 1.427 ;
      RECT 1.227 0.681 1.277 0.903 ;
      RECT 1.039 0.953 1.089 1.213 ;
      RECT 0.583 1.213 1.089 1.263 ;
      RECT 0.735 0.098 1.089 0.148 ;
      RECT 0.735 0.148 0.785 0.501 ;
      RECT 1.039 0.148 1.089 0.431 ;
      RECT 0.279 0.598 0.937 0.648 ;
      RECT 0.583 0.181 0.633 0.598 ;
      RECT 0.887 0.208 0.937 0.598 ;
      RECT 0.279 0.178 0.329 0.598 ;
    LAYER PO ;
      RECT 1.125 0.101 1.155 1.469 ;
      RECT 1.885 0.101 1.915 1.469 ;
      RECT 0.517 0.101 0.547 1.567 ;
      RECT 1.581 0.069 1.611 1.608 ;
      RECT 0.821 0.101 0.851 1.469 ;
      RECT 0.669 0.101 0.699 1.469 ;
      RECT 0.213 0.101 0.243 1.469 ;
      RECT 0.365 0.101 0.395 1.469 ;
      RECT 1.277 0.101 1.307 1.469 ;
      RECT 1.733 0.101 1.763 1.469 ;
      RECT 1.429 0.069 1.459 1.608 ;
      RECT 0.973 0.101 1.003 1.469 ;
      RECT 0.061 0.101 0.091 1.469 ;
    LAYER CO ;
      RECT 0.587 1.23 0.629 1.272 ;
      RECT 0.587 1.322 0.629 1.364 ;
      RECT 0.587 0.423 0.629 0.465 ;
      RECT 0.739 0.239 0.781 0.281 ;
      RECT 1.423 0.635 1.465 0.677 ;
      RECT 0.587 0.331 0.629 0.373 ;
      RECT 1.575 0.635 1.617 0.677 ;
      RECT 0.587 1.138 0.629 1.18 ;
      RECT 1.195 0.362 1.237 0.404 ;
      RECT 1.195 1.355 1.237 1.397 ;
      RECT 0.587 0.239 0.629 0.281 ;
      RECT 0.739 0.423 0.781 0.465 ;
      RECT 0.891 0.239 0.933 0.281 ;
      RECT 0.283 0.239 0.325 0.281 ;
      RECT 0.739 0.331 0.781 0.373 ;
      RECT 1.195 1.263 1.237 1.305 ;
      RECT 1.043 0.178 1.085 0.22 ;
      RECT 0.891 0.331 0.933 0.373 ;
      RECT 1.195 0.27 1.237 0.312 ;
      RECT 1.043 0.27 1.085 0.312 ;
      RECT 0.283 0.423 0.325 0.465 ;
      RECT 0.891 0.423 0.933 0.465 ;
      RECT 1.043 0.362 1.085 0.404 ;
      RECT 0.283 0.331 0.325 0.373 ;
    LAYER NWELL ;
      RECT -0.135 0.679 2.092 1.787 ;
  END
END OA221X2_RVT

MACRO NAND4X1_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1.824 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 1.043 0.857 1.085 ;
      LAYER M1 ;
        RECT 0.705 1.089 0.815 1.119 ;
        RECT 0.705 1.039 0.877 1.089 ;
        RECT 0.705 1.009 0.815 1.039 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0183 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.738 0.705 0.78 ;
      LAYER M1 ;
        RECT 0.553 0.785 0.663 0.815 ;
        RECT 0.553 0.735 0.725 0.785 ;
        RECT 0.553 0.705 0.663 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0183 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 1.043 0.553 1.085 ;
      LAYER M1 ;
        RECT 0.401 1.089 0.511 1.119 ;
        RECT 0.401 1.039 0.573 1.089 ;
        RECT 0.401 1.009 0.511 1.039 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0183 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.738 0.401 0.78 ;
      LAYER M1 ;
        RECT 0.249 0.785 0.359 0.815 ;
        RECT 0.249 0.735 0.421 0.785 ;
        RECT 0.249 0.705 0.359 0.735 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0183 ;
  END A4
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.347 0.15 1.389 0.192 ;
        RECT 1.347 0.242 1.389 0.284 ;
        RECT 1.347 0.334 1.389 0.376 ;
        RECT 1.347 0.426 1.389 0.468 ;
        RECT 1.347 0.936 1.389 0.978 ;
        RECT 1.347 1.028 1.389 1.07 ;
        RECT 1.347 1.12 1.389 1.162 ;
        RECT 1.347 1.212 1.389 1.254 ;
        RECT 1.347 1.304 1.389 1.346 ;
        RECT 1.347 1.396 1.389 1.438 ;
        RECT 1.347 1.488 1.389 1.53 ;
      LAYER M1 ;
        RECT 1.343 0.876 1.393 1.565 ;
        RECT 1.343 0.826 1.64 0.876 ;
        RECT 1.59 0.815 1.64 0.826 ;
        RECT 1.59 0.705 1.727 0.815 ;
        RECT 1.59 0.564 1.64 0.705 ;
        RECT 1.343 0.514 1.64 0.564 ;
        RECT 1.343 0.115 1.393 0.514 ;
    END
    ANTENNADIFFAREA 0.1244 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 1.499 1.028 1.541 1.07 ;
        RECT 1.499 1.12 1.541 1.162 ;
        RECT 1.043 1.203 1.085 1.245 ;
        RECT 1.499 1.212 1.541 1.254 ;
        RECT 1.043 1.295 1.085 1.337 ;
        RECT 1.499 1.304 1.541 1.346 ;
        RECT 1.043 1.387 1.085 1.429 ;
        RECT 1.499 1.396 1.541 1.438 ;
        RECT 0.435 1.397 0.477 1.439 ;
        RECT 0.739 1.397 0.781 1.439 ;
        RECT 1.043 1.479 1.085 1.521 ;
        RECT 1.499 1.488 1.541 1.53 ;
        RECT 0.435 1.489 0.477 1.531 ;
        RECT 0.739 1.489 0.781 1.531 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 1.824 1.702 ;
        RECT 0.431 1.377 0.481 1.642 ;
        RECT 0.735 1.377 0.785 1.642 ;
        RECT 1.039 1.183 1.089 1.642 ;
        RECT 1.495 1.008 1.545 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 0.283 0.141 0.325 0.183 ;
        RECT 1.043 0.142 1.085 0.184 ;
        RECT 1.499 0.152 1.541 0.194 ;
        RECT 0.283 0.233 0.325 0.275 ;
        RECT 1.043 0.234 1.085 0.276 ;
        RECT 1.499 0.244 1.541 0.286 ;
        RECT 0.283 0.325 0.325 0.367 ;
        RECT 1.499 0.336 1.541 0.378 ;
        RECT 0.283 0.417 0.325 0.459 ;
      LAYER M1 ;
        RECT 0.279 0.03 0.329 0.479 ;
        RECT 1.495 0.03 1.545 0.413 ;
        RECT 1.039 0.03 1.089 0.296 ;
        RECT 0 -0.03 1.824 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 0.587 1.489 0.629 1.531 ;
      RECT 0.283 1.489 0.325 1.531 ;
      RECT 1.195 0.142 1.237 0.184 ;
      RECT 0.891 0.233 0.933 0.275 ;
      RECT 0.891 1.489 0.933 1.531 ;
      RECT 1.423 0.618 1.465 0.66 ;
      RECT 0.891 0.141 0.933 0.183 ;
      RECT 1.119 0.741 1.161 0.783 ;
      RECT 1.195 1.295 1.237 1.337 ;
      RECT 1.195 1.479 1.237 1.521 ;
      RECT 1.195 1.203 1.237 1.245 ;
      RECT 1.195 1.295 1.237 1.337 ;
      RECT 1.195 1.387 1.237 1.429 ;
      RECT 1.195 1.203 1.237 1.245 ;
      RECT 1.195 1.387 1.237 1.429 ;
      RECT 1.195 1.479 1.237 1.521 ;
      RECT 0.891 0.325 0.933 0.367 ;
      RECT 0.891 0.417 0.933 0.459 ;
      RECT 0.891 1.397 0.933 1.439 ;
      RECT 0.587 1.397 0.629 1.439 ;
      RECT 0.283 1.397 0.325 1.439 ;
      RECT 1.195 0.142 1.237 0.184 ;
      RECT 1.195 0.234 1.237 0.276 ;
    LAYER M1 ;
      RECT 0.927 0.737 1.181 0.787 ;
      RECT 0.279 1.327 0.329 1.551 ;
      RECT 0.583 1.327 0.633 1.551 ;
      RECT 0.279 1.277 0.977 1.327 ;
      RECT 0.887 0.587 0.977 0.637 ;
      RECT 0.887 1.327 0.937 1.551 ;
      RECT 0.887 0.121 0.937 0.587 ;
      RECT 0.927 0.787 0.977 1.277 ;
      RECT 0.927 0.637 0.977 0.737 ;
      RECT 1.231 0.614 1.485 0.664 ;
      RECT 1.191 0.906 1.241 1.556 ;
      RECT 1.191 0.856 1.281 0.906 ;
      RECT 1.191 0.114 1.241 0.455 ;
      RECT 1.191 0.455 1.281 0.505 ;
      RECT 1.231 0.664 1.281 0.856 ;
      RECT 1.231 0.505 1.281 0.614 ;
    LAYER PO ;
      RECT 0.365 0.071 0.395 1.61 ;
      RECT 0.517 0.071 0.547 1.61 ;
      RECT 0.669 0.071 0.699 1.61 ;
      RECT 0.213 0.071 0.243 1.61 ;
      RECT 1.277 0.064 1.307 1.6 ;
      RECT 1.125 0.064 1.155 1.61 ;
      RECT 0.821 0.071 0.851 1.61 ;
      RECT 1.581 0.071 1.611 1.61 ;
      RECT 0.061 0.071 0.091 1.61 ;
      RECT 1.429 0.072 1.459 1.61 ;
      RECT 0.973 0.071 1.003 1.61 ;
      RECT 1.733 0.064 1.763 1.6 ;
    LAYER NWELL ;
      RECT -0.115 0.679 1.959 1.773 ;
  END
END NAND4X1_RVT

MACRO OR4X4_RVT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2.584 BY 1.672 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.359 0.548 0.401 0.59 ;
      LAYER M1 ;
        RECT 0.249 0.528 0.417 0.663 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0315 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.511 0.548 0.553 0.59 ;
      LAYER M1 ;
        RECT 0.401 0.857 0.557 0.967 ;
        RECT 0.507 0.528 0.557 0.857 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0315 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.663 0.548 0.705 0.59 ;
      LAYER M1 ;
        RECT 0.657 0.705 0.815 0.815 ;
        RECT 0.659 0.528 0.709 0.705 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0315 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 0.815 0.548 0.857 0.59 ;
      LAYER M1 ;
        RECT 0.811 0.511 0.861 0.61 ;
        RECT 0.807 0.4 0.967 0.511 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0315 ;
  END A4
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER CO ;
        RECT 1.803 0.151 1.845 0.193 ;
        RECT 2.107 0.151 2.149 0.193 ;
        RECT 1.803 0.245 1.845 0.287 ;
        RECT 2.107 0.245 2.149 0.287 ;
        RECT 1.803 0.337 1.845 0.379 ;
        RECT 2.107 0.337 2.149 0.379 ;
        RECT 1.803 0.43 1.845 0.472 ;
        RECT 2.107 0.43 2.149 0.472 ;
        RECT 1.803 0.915 1.845 0.957 ;
        RECT 2.107 0.915 2.149 0.957 ;
        RECT 1.803 1.009 1.845 1.051 ;
        RECT 2.107 1.009 2.149 1.051 ;
        RECT 1.803 1.101 1.845 1.143 ;
        RECT 2.107 1.101 2.149 1.143 ;
        RECT 1.803 1.194 1.845 1.236 ;
        RECT 2.107 1.194 2.149 1.236 ;
        RECT 1.803 1.286 1.845 1.328 ;
        RECT 2.107 1.286 2.149 1.328 ;
        RECT 1.803 1.38 1.845 1.422 ;
        RECT 2.107 1.38 2.149 1.422 ;
        RECT 1.803 1.472 1.845 1.514 ;
        RECT 2.107 1.472 2.149 1.514 ;
      LAYER M1 ;
        RECT 1.799 0.945 1.849 1.534 ;
        RECT 2.103 0.945 2.153 1.534 ;
        RECT 1.799 0.895 2.439 0.945 ;
        RECT 2.389 0.49 2.439 0.895 ;
        RECT 1.799 0.49 1.849 0.492 ;
        RECT 2.103 0.49 2.153 0.492 ;
        RECT 1.799 0.44 2.439 0.49 ;
        RECT 1.799 0.131 1.849 0.44 ;
        RECT 2.103 0.131 2.153 0.44 ;
        RECT 2.389 0.359 2.439 0.44 ;
        RECT 2.377 0.249 2.487 0.359 ;
    END
    ANTENNADIFFAREA 0.2976 ;
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER CO ;
        RECT 0.283 0.744 0.325 0.786 ;
        RECT 0.283 0.838 0.325 0.88 ;
        RECT 1.043 0.901 1.085 0.943 ;
        RECT 0.283 0.93 0.325 0.972 ;
        RECT 1.043 0.993 1.085 1.035 ;
        RECT 0.283 1.024 0.325 1.066 ;
        RECT 1.347 1.025 1.389 1.067 ;
        RECT 1.043 1.085 1.085 1.127 ;
        RECT 2.259 1.115 2.301 1.157 ;
        RECT 0.283 1.116 0.325 1.158 ;
        RECT 1.651 1.116 1.693 1.158 ;
        RECT 1.955 1.116 1.997 1.158 ;
        RECT 1.347 1.117 1.389 1.159 ;
        RECT 2.259 1.208 2.301 1.25 ;
        RECT 0.283 1.209 0.325 1.251 ;
        RECT 1.347 1.209 1.389 1.251 ;
        RECT 1.651 1.209 1.693 1.251 ;
        RECT 1.955 1.209 1.997 1.251 ;
        RECT 2.259 1.3 2.301 1.342 ;
        RECT 0.283 1.301 0.325 1.343 ;
        RECT 1.347 1.301 1.389 1.343 ;
        RECT 1.651 1.301 1.693 1.343 ;
        RECT 1.955 1.301 1.997 1.343 ;
        RECT 2.259 1.394 2.301 1.436 ;
        RECT 0.283 1.395 0.325 1.437 ;
        RECT 1.347 1.395 1.389 1.437 ;
        RECT 1.651 1.395 1.693 1.437 ;
        RECT 1.955 1.395 1.997 1.437 ;
        RECT 2.259 1.486 2.301 1.528 ;
        RECT 0.283 1.487 0.325 1.529 ;
        RECT 1.347 1.487 1.389 1.529 ;
        RECT 1.651 1.487 1.693 1.529 ;
        RECT 1.955 1.487 1.997 1.529 ;
        RECT 0.055 1.651 0.097 1.693 ;
        RECT 0.207 1.651 0.249 1.693 ;
        RECT 0.359 1.651 0.401 1.693 ;
        RECT 0.511 1.651 0.553 1.693 ;
        RECT 0.663 1.651 0.705 1.693 ;
        RECT 0.815 1.651 0.857 1.693 ;
        RECT 0.967 1.651 1.009 1.693 ;
        RECT 1.119 1.651 1.161 1.693 ;
        RECT 1.271 1.651 1.313 1.693 ;
        RECT 1.423 1.651 1.465 1.693 ;
        RECT 1.575 1.651 1.617 1.693 ;
        RECT 1.727 1.651 1.769 1.693 ;
        RECT 1.879 1.651 1.921 1.693 ;
        RECT 2.031 1.651 2.073 1.693 ;
        RECT 2.183 1.651 2.225 1.693 ;
        RECT 2.335 1.651 2.377 1.693 ;
        RECT 2.487 1.651 2.529 1.693 ;
      LAYER M1 ;
        RECT 0 1.642 2.584 1.702 ;
        RECT 0.279 0.724 0.329 1.642 ;
        RECT 1.039 0.881 1.089 1.642 ;
        RECT 1.343 1.005 1.393 1.642 ;
        RECT 1.647 1.096 1.697 1.642 ;
        RECT 1.951 1.096 2.001 1.642 ;
        RECT 2.255 1.095 2.305 1.642 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER CO ;
        RECT 0.055 -0.021 0.097 0.021 ;
        RECT 0.207 -0.021 0.249 0.021 ;
        RECT 0.359 -0.021 0.401 0.021 ;
        RECT 0.511 -0.021 0.553 0.021 ;
        RECT 0.663 -0.021 0.705 0.021 ;
        RECT 0.815 -0.021 0.857 0.021 ;
        RECT 0.967 -0.021 1.009 0.021 ;
        RECT 1.119 -0.021 1.161 0.021 ;
        RECT 1.271 -0.021 1.313 0.021 ;
        RECT 1.423 -0.021 1.465 0.021 ;
        RECT 1.575 -0.021 1.617 0.021 ;
        RECT 1.727 -0.021 1.769 0.021 ;
        RECT 1.879 -0.021 1.921 0.021 ;
        RECT 2.031 -0.021 2.073 0.021 ;
        RECT 2.183 -0.021 2.225 0.021 ;
        RECT 2.335 -0.021 2.377 0.021 ;
        RECT 2.487 -0.021 2.529 0.021 ;
        RECT 0.435 0.138 0.477 0.18 ;
        RECT 0.739 0.138 0.781 0.18 ;
        RECT 1.043 0.141 1.085 0.183 ;
        RECT 2.259 0.164 2.301 0.206 ;
        RECT 1.347 0.165 1.389 0.207 ;
        RECT 1.651 0.165 1.693 0.207 ;
        RECT 1.955 0.165 1.997 0.207 ;
        RECT 2.259 0.256 2.301 0.298 ;
        RECT 1.347 0.257 1.389 0.299 ;
        RECT 1.651 0.257 1.693 0.299 ;
        RECT 1.955 0.257 1.997 0.299 ;
      LAYER M1 ;
        RECT 1.343 0.03 1.393 0.319 ;
        RECT 1.647 0.03 1.697 0.319 ;
        RECT 1.951 0.03 2.001 0.319 ;
        RECT 2.255 0.03 2.305 0.318 ;
        RECT 1.039 0.03 1.089 0.203 ;
        RECT 0.431 0.03 0.481 0.2 ;
        RECT 0.735 0.03 0.785 0.2 ;
        RECT 0 -0.03 2.584 0.03 ;
    END
  END VSS
  OBS
    LAYER CO ;
      RECT 2.031 0.67 2.073 0.712 ;
      RECT 1.119 0.67 1.161 0.712 ;
      RECT 1.195 0.245 1.237 0.287 ;
      RECT 1.195 0.151 1.237 0.193 ;
      RECT 1.195 0.989 1.237 1.031 ;
      RECT 1.195 0.897 1.237 0.939 ;
      RECT 1.195 0.803 1.237 0.845 ;
      RECT 1.879 0.67 1.921 0.712 ;
      RECT 1.499 0.334 1.541 0.376 ;
      RECT 1.499 0.242 1.541 0.284 ;
      RECT 1.499 0.148 1.541 0.19 ;
      RECT 2.183 0.67 2.225 0.712 ;
      RECT 1.499 0.427 1.541 0.469 ;
      RECT 1.499 1.458 1.541 1.5 ;
      RECT 1.499 1.366 1.541 1.408 ;
      RECT 1.423 0.667 1.465 0.709 ;
      RECT 1.499 1.272 1.541 1.314 ;
      RECT 1.499 1.18 1.541 1.222 ;
      RECT 1.499 1.087 1.541 1.129 ;
      RECT 1.499 0.995 1.541 1.037 ;
      RECT 1.727 0.67 1.769 0.712 ;
      RECT 1.499 0.901 1.541 0.943 ;
      RECT 0.891 0.189 0.933 0.231 ;
      RECT 0.283 0.189 0.325 0.231 ;
      RECT 0.891 1.458 0.933 1.5 ;
      RECT 0.891 1.366 0.933 1.408 ;
      RECT 0.891 1.272 0.933 1.314 ;
      RECT 0.891 1.18 0.933 1.222 ;
      RECT 0.891 1.087 0.933 1.129 ;
      RECT 0.587 0.189 0.629 0.231 ;
      RECT 0.891 0.995 0.933 1.037 ;
      RECT 0.891 0.903 0.933 0.945 ;
      RECT 0.891 0.811 0.933 0.853 ;
    LAYER M1 ;
      RECT 1.618 0.666 2.245 0.716 ;
      RECT 1.495 0.556 1.545 0.557 ;
      RECT 1.495 0.128 1.545 0.506 ;
      RECT 1.495 0.947 1.545 1.535 ;
      RECT 1.495 0.881 1.545 0.897 ;
      RECT 1.495 0.897 1.668 0.947 ;
      RECT 1.618 0.716 1.668 0.897 ;
      RECT 1.495 0.506 1.668 0.556 ;
      RECT 1.618 0.556 1.668 0.666 ;
      RECT 1.029 0.666 1.181 0.716 ;
      RECT 1.029 0.303 1.079 0.666 ;
      RECT 0.279 0.253 1.079 0.303 ;
      RECT 1.029 0.716 1.079 0.731 ;
      RECT 0.887 0.731 1.079 0.781 ;
      RECT 0.279 0.169 0.329 0.253 ;
      RECT 0.583 0.169 0.633 0.253 ;
      RECT 0.887 0.168 0.937 0.253 ;
      RECT 0.887 0.781 0.937 1.535 ;
      RECT 1.34 0.663 1.485 0.713 ;
      RECT 1.34 0.477 1.39 0.663 ;
      RECT 1.192 0.452 1.39 0.477 ;
      RECT 1.191 0.427 1.39 0.452 ;
      RECT 1.34 0.713 1.39 0.803 ;
      RECT 1.191 0.803 1.39 0.853 ;
      RECT 1.191 0.853 1.241 1.051 ;
      RECT 1.191 0.783 1.241 0.803 ;
      RECT 1.191 0.131 1.241 0.427 ;
    LAYER PO ;
      RECT 2.037 0.071 2.067 1.612 ;
      RECT 1.885 0.071 1.915 1.612 ;
      RECT 1.733 0.071 1.763 1.612 ;
      RECT 2.189 0.071 2.219 1.612 ;
      RECT 2.341 0.071 2.371 1.612 ;
      RECT 1.581 0.071 1.611 1.612 ;
      RECT 1.125 0.071 1.155 1.612 ;
      RECT 1.277 0.071 1.307 1.612 ;
      RECT 1.429 0.071 1.459 1.61 ;
      RECT 0.973 0.061 1.003 1.61 ;
      RECT 0.061 0.061 0.091 1.61 ;
      RECT 2.493 0.072 2.523 1.61 ;
      RECT 0.821 0.061 0.851 1.61 ;
      RECT 0.213 0.061 0.243 1.61 ;
      RECT 0.669 0.061 0.699 1.61 ;
      RECT 0.365 0.061 0.395 1.61 ;
      RECT 0.517 0.061 0.547 1.61 ;
    LAYER NWELL ;
      RECT -0.115 0.679 2.699 1.801 ;
      RECT 0.198 0.565 1.018 0.679 ;
  END
END OR4X4_RVT

END LIBRARY
